<!DOCTYPE html><html><head><meta charset="UTF-8"><title>Spice-Up - WebViewer</title><meta name="viewport" content="width=device-width, initial-scale=1"/></head><style>.slides{background-color: #363B3E;}html, body{background-color: #363B3E;}#content{display: none;}.slide{ background-color: lightgray; position: relative; overflow: hidden; margin-bottom: 16px; margin-left: auto; margin-right: auto; border: solid 1px #0E0F10; border-radius: 12px;}.slide-16-9{min-width: 1920px; max-width: 1920px; min-height: 1080px; max-height: 1080px;}.slide-16-10{min-width: 1920px; max-width: 1920px; min-height: 1200px; max-height: 1200px;}.slide-4-3{min-width: 1920px; max-width: 1920px; min-height: 1440px; max-height: 1440px;}.slide-3-2{min-width: 1920px; max-width: 1920px; min-height: 1280px; max-height: 1280px;}.slide-5-4{min-width: 1920px; max-width: 1920px; min-height: 1536px; max-height: 1536px;}.canvas-item{position: absolute; display: flex;}text-item{white-space: pre-wrap;}text-item span{align-self: center;}</style><script>if (!String.build){String.build=function (format){var args=Array.prototype.slice.call (arguments, 1); return format.replace (/{(\d+)}/g, function (match, number){return typeof args[number] !='undefined' ? args[number] : match;});};}function base64Decode(str){return decodeURIComponent(Array.prototype.map.call(atob(str), function(c){return '%' + ('00' + c.charCodeAt(0).toString(16)).slice(-2);}).join(''));}function makeIdEditable (id){get (id).contentEditable="true";}function get (id){return document.getElementById(id);}function downloadString (element, fileName, mime){var dlAnchorElem=document.getElementById ('download-anchor'); if (dlAnchorElem===null){document.getElementById ("body").innerHTML +='<a id="download-anchor" style="display:none"></a>'; dlAnchorElem=document.getElementById ('download-anchor');}var dataStr="data:" + mime + ";charset=utf-8," + encodeURIComponent(element); var dlAnchorElem=document.getElementById ('download-anchor'); dlAnchorElem.setAttribute ("href", dataStr); dlAnchorElem.setAttribute ("download", fileName); dlAnchorElem.click ();}</script><body id="body"> <h1 style="color: #dfdfdf; font-family: sans-serif; text-align: center; width: 100%; margin-top: 200px; font-size: 3em"> Loading presentation... </h1> <content id="content">
{"current-slide":1, "preview-slide":0, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(360deg, #606c88 0%, #3f4c6b 49%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/45-degree-fabric-dark.png" , "transition": 0, "items": [{"x": -638,"y": 73,"w": 2767,"h": 472,"type":"text","text": "","text-data": "RmluYWwgUHJvamVjdA==","font": "raleway","color": "#ffffff","font-size": 42, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -648,"y": 902,"w": 2784,"h": 315,"type":"text","text": "","text-data": "w4FsdmFybyBHYWxpc3Rlbw==","font": "raleway","color": "#fff394","font-size": 28, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -638,"y": 409,"w": 2769,"h": 190,"type":"text","text": "","text-data": "QWR2YW5jZWQgQ29tcHV0ZXIgQXJjaGl0ZWN0dXJl","font": "raleway","color": "#ffffff","font-size": 21, "font-style":"regular", "justification": 1, "align": 1 }
,{"x": -641,"y": 1105,"w": 2774,"h": 334,"type":"text","text": "","text-data": "QmFjaGVsb3IgZGVncmVlIGluIGNvbXB1dGVyIGVuZ2luZWVyaW5nClRVIFdpZW4gRXJhc211cyAxOS8yMA==","font": "raleway","color": "#ffffff","font-size": 16, "font-style":"regular", "justification": 1, "align": 1 }
], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nJx9d5xlRZX/t+57Pd09OTADDMwAg2SGIJIzA4gEEUTWVRQjrhhYdXXN66qoqGta8ypGVDCAICgoiIAokkGGMENmYAYmhw7T3bd+f1Sdc76n7m3083s6vNc3VJ3vyXWqbt1wwGEnXt7pmbgIQAAQUUegCsif/CMCMQIxRABAxafqgBhiOpYOBgTEWCOEChFRm7ZGQ/4rAhEIVbo5xlrbDSGkPgFpIwYg5DsCEGMIIcR0TQwBIcZ8H9K9EYjpb2R6QogxpibgMEbEGBACncg/Y/0PcAckniGEEJDp8ezLaB1uACFUueuYz0KgteGGkC+4mavSltwWQ2qPcCM1HIywOkZU0OaZ1nHlXWcZVQFADCIrweB524Y7qGxFNxg3X6dcLHETnxNuAJkh0mKMYwihE5JOKW6mKxhvIx3OHKwKGcY6pOPGv4Sridfdl48HBEDpJj5kXmfcooRZ3ElsSbej6oHwPOt55K4Sf6rnwR2EusA2iACgdrizQGJADHFsbPi6bqenf1Ho9E7U9ioAqIFQqdKiuJ8/CVXFf2XmCDv5SkWUrgkddzxkBUrtkbIwCY4coscsCsgKpcLMjgtiYLE2BXU00bESe9tHDLQjlEUSRdlGaO+X+IHnxW2GlXAnow3OY+gVAOrMh0RjiBFiaMgaiA71nZVZFDe0yBoAUAGh6pBjF4dQUmz3pn7zzaS/wfG82QIrdxWyybXhFnrFuctdIV8veOVbeQ53reMPnYzCR24jtuEu+KX4zJZCFcllZ/0JwbwATNYetzhHZB/tnWWMYzDHS7wVOkLQWAJqw4XMCu6jehACOqNhUTcZLEwuHGQg0U3aC57ZQWKGv8e355mfDCb9TwQrXFDH4xwia0VFv6PLROyw+OhScNJX7ruqgMzgRjcS9aIxi9v2mORG359FHcNNf9ht0v3z4s6GEBKOGEk5udsIRNSeT2W2FgS3NC3hODgaLUtzB3Kw4SwCDohG/Xy9yiECKQhBFdU5pcAMYdzSffTnHbtj5knWqUA6EZEwl86bronZsY6HO+mqKrS1E7OD5/40UyTqiSZzFEJrS1Bm3LXcK7jlPpieCk2qFqFoJ9KfrLuaW+Qcy+Ng2YQQ0NUsJgsrhI562BTlrS9RWBO1MTBdT0yVoQwbNMwTGvXJa8uwxStKZpR40hBJaMQMERozpujDhMKRgYQQOg5boOaDOjJS2iC8ENwZpxpUEXlDQbO0ITx2H6GX8WRFYafscOf+lD0lbu/kmffeQdGtKpeQnVDGTIqfOqxacKeGQtk2ooRL6pYcLstbrnd4x8MtMpFoXSWZ5L5UgE4XA2KWofmhbAPSLmp3veHO7bnAUcqasUfPD+cgmT8KlngDczh8mWDUgJbtsHRCJe5KeOfloMPiAAsooVIdr1K2rlZh0VCMovDgFlkKaNG8cxrn53/6d6TzPiJpRItjpgixLvoOvn3rODPDMgfP0aJPSv18NMPzYItArMkPMztqOhYzbYI1FnwRrZVoUNtxVWbmTRlp23DLdXkIU2ZBTmGyZqhTTpE/4nlkKvgNcL6eIrjDLfyQf4KPjEL+dn1yEGhxFKDTgfgTOhl3hUafkkWWhpfvj0ob98/66B1VjIxb7CPhjdm4Ghlki/247KfxIQx8TPps6HFlt0FkJcP/MjAYL1wwU5WpE1eil4Xg7jpmEY119NE1AeQagyioGYVWKMrxIR9zvwM0W1AlZpDwSsaRj9ulg77YBvO0yncxVBaKKa/e6Tx6x+7VqCaKgiYuTXvFWxc80BS0hU8ocZeAS9zpvC/6BcRy7K24M152WBEet3NezX5jnWsvGn0Yd0U8MvI1g9UMQCJ+ca2Ttx4sjpkusCtNw2JfZHZOsNTzegwpi8z01GMkdwc6Yxgfd1B6zDhdQyXu8qMOZBzcKg/GTTruGFHg1mPZ+Stu4UM9Pm51hBHdJtUBkl7b3QGoOtkJBWrPlKoxvGBP4yK/nI/FtW2f4PkepMIPOk5eMBRRIafRbjxXtu+iTlGQDQG5ellgKbw7RSWX0geYQykdQkDzehvQ/gPchfEUuHWIyAGixK0k0zSW4mZZOmbn7tpwBz0nRWXjEaBFO8efHHDYUJxIgkBqxw14eaNCdHrG1zIzhN7o2VPRX42sJ+N2WQHhrqp8i2RWgnU83BIwKuubnH0Dt8hKayuSyQGxqOX5mlURdLJ+OXlXnXGuF3o6iAC6CFWeXqTpyzbPp7eX0SqTESpwrcMMORPZcAq+9Cr3IyB7Oone4o0t8lt0yAaeo6qJPzFAZBVpmCV027iSpy/LT0uEYNyhwB3La00p9W8ZQ2tUqOw+dbDPh5uiCxcTBX3VyVGjMllJu7HOgo8IoZtxc20l0D9xBoSHs8GC93KNZnWa2Uiw8bWTdJ+wxTCxg/TDH7rGZU1krIkiz8/Ma3Nw4swYHxl/eTzKDJ30XRE/GXc+5grV9LfwCgAiDYXlo/e34YZzFEZzQKhkFqcqeC+sItycYTt5S/9Rg2wZ5AKqWMUxHms1PbcRbYIPbHxZ0I7gcZ2NKYpXxhwZxVGVY3dHGyDjRzkvyurqA/UYZDzulF3H4akG4RlY4HbjbzKk8XCP+2GhcHu14bZOC9wMm6+VMTfXPYwHbMAJQg3lM4CoMyIWbXy/pfNg+DlbKHG7sS7gMk43FBwPN/XtDLHOjo70wmUU1p7T42htR5K7BXnCVuIOpUGb3geZAi6d6D/AHeuxQpfJDmLxrTTntpXPrJOG1+Nm2yA9Z7NSfawd7iBZBs3yiJOrUhY4lp21Eeo9rPBAorDQEu0fCcScinhZYT4c8+03p6zkHVlRjeVAqMxhNVJyabucdTG6FJ8r4I2Hm6OS4GwTKrfPGCuIoulaAC1WKWNbeEJ487ekg45Opk3XaVB7yjPpU5SjLOS14S6UOSal8wpKPJY1HSUdPMTgPqjAHFg/nEOFtif9JhFz6v0PcEeSG9CCmz+yaMxkmsiuwQ7H6SkZVaNG1Ya76E+vcbocYMsacn9BsMqnxC0kx+xfWKeRF9QJLaIz3hnaVLcEnYQ7BARdZ2HjrUCEmTAdAzTdYcDmgSQ7aEzhKBYBIdGpdCSAr9iYV0++h+smwch01wkWZiQVHitKyzTlQituyx4SnuBmXoSeCBs6UPGSg5ziFt7RFJYqlBe84ZFJK0qD9aIKsvjUT10Sj7JihxC9EjkZRuE2uY58PA8jQmzBLddFpgFJB9QpEn/4flFs5kOQWQx1JVkdcvtydaiANtysozHmehs7hnbDlUzJrzoeR89j0Y8aJ4AyqyhwK42cNeSA2ghr0g+RnepCcr4MlnZtKHG7jN0wmY6VjhyQgm2MMVYxjpF3NE8VNHpzhJEvOS/TdelE8jcp1QowRTcscTw5gaNXYjKnW6l1XWEHdyo7HfOMrq7iLrRhiqx406xHM4CMO/AaAWFkUOZxBEm4LQ0MukaCcbNhRjUGR5dGfY4AUNyu4EW8pPhPBLcMbWSYAo9Z8UjqGYr7QoWQdSOlqXI2JtyxmDljGjxRDrdzWjwMjYQbVo/yOmg/fRcUSSHrhCIsEDb1XPS/XPbtdLykO0feUBhyEkZd6GCTNbac4B/gdgV14gLXsaQ9yjgtO4rwGSfrL9kMOYoQOmTbIbdXhW4IVfBjT1Eo8Y55kiVGaKVZCM1M0dVfta0MbIy3lJkRtoiHGVz6VJjHBbToae1KATSaV+c55+ylJROR5owjlRMQNE21dtv8WsI9hjpmrxuCpXcyfuaLteJdA7HELQL1mQxH+ViPZdxjmS6Ti7JJQ3M03JnH5lvEkXVM2RFg60egDsamXYPeF5FoiA43OSFxeDyMoGHl+HUdwk2GkfAKbhaTzUYYbssKNIvI3kuoV9zSJ+EyPbIoz9Pvkin5JeWJVnN49rcOv8kYk+FF42sDN6i9gBhH8zfT21x4mHDVlD3B2mW+UPsJpthS8PyiTCTGWh+hiDFpFORpFe3AKUk041NvY1NIgSKUVd9Z6SV65/uco6CiZKsiyUf6kvb8HL5+iiKPjVFpCa5Lr3hWRJKA2nAj4666ieaqo8YflI6Mm8au2loAefU23HU7bpcOkpKysnBay4VYjhItuLVlqhHo0nuOrqFKY2bNOJMRPC9urslwNBNnzvLWnICcnyMQzahe6CnjZswQnRXHpkaAgla0y5t1PRu/mzFk/pmQzEaU7gK31gzgMQHwK0WznVg0IEcq2ETWZPAwWedfhYOWekzCHYinIS9u4+eyDEuSf5U56gWhFyErTGrcFbScQiREzWWuBWNIoQWUt/byWj5mBS5mjDEq+HvHmWGIrByhYGYDdyDcgRhr16X4xtlTGw887sb4lXHHEneF6IwrEpyWuowrtvqIou1rBJVugtKkUZFxCy0qc8KtfQW9rImb8QS6poVXwa6zbMrPCo0r78aYvGVKnO/Vir+fvXA5pV5jzsGtCs3ZjVN9DlqEB+PaB10DjI9brxPZCe78W7OdcYKQXKNDr0p5FmlU4OlRrLGKKewSSG67YBpADiEAAqphCHJIvOoYonM2osg8DZuPB+/d6CTRVCiKa1MYEjxdLFxpp3EOxT2C2xuwTjuKUELGnTFwNOHZg3bc9q3j57aPU3JRmJwRuIVATYPxvBQlbJNZbW1o5kH80eEWDTn0IpslasctPCrwadYZPN+Z5nKmZDzcPNxtw936W3BTX+40BSfG7XRHMJOeuxpAm1McT9ZtuEHt8ZA3EC8YF+tW6TQoaOi5slZluOxahG4IIWilX05wxCk6ST5GvDhHCll0IgKTTIOmgAA9FutRaHGVGaVj6OBnLKwBmKEI0CxQFkDMBqm+gY2V6G3LQFyKScx2uGGr9oqUVlLWoFEFlhrWY0AcQ3T1FWTcocBt0aIZhIupQ+kreuV06y0UW+EQ4/PgjjADkXYrvs7uN3lbcSxIRtg6S1NkHbpwqzR0+jh9sdkt7Vd2aShw29g999lYQSwNFXzhLLDiSEvfqv8cCHJQqaMtCnS4haeMoQ13hOq40IvgFvfpkgYALquJ0ePmNl12S7IuAiNUl6vYtcxCPHzuMFKj7E358WbNKiR9IkYosCYBOqVaesKCSL+6MJLXj8gVRmujqsCyNoGVXhfqEMXQbdWfME3oI5zsRAGkBTGZ4W7eHoVHJ4Nuw63LfC0a+GGP4C5pIwNnZZPaREvWlKrshWNwuCPRHsbHk5XUfo/jbNiR8hqa8lNmNnJ/qDx9doM5L+eoYlO3YjFrEKp8m7RLfZZZQzlcUxYUAabAbSgpWmtwK3GM054LbqHgpdElQ6LGStwW3I72hj7na90w1WwbMYYuEIM8huyMPMTcHnmhUHKtxTvJYVYoO9AcQyrDYIbrIgItC45yacjkiEeN1H2E1SLqZj/y0EzMy3gjyPNnxgNmVC57Ytq5Mk3Rn+lwuGvXun5I2fmJPytSpWP86LE6QsEdkbFWisvRDkBXQObMTessGmHYubC8GxpO1wfI3mUEKClmPZZ1tibjDP6eQFUPKZijnAGQ/ux6w22ORO9BQXMIaSMYNUhb2+EXOJV6zo6yBZ+jj+6XoRgkqhPPFHf6OyjuwnETbt3cRofVMKfacAgALyUvcY/nq4lZ3rmRnCPybEhzj4l0sZ9nLiJV5JWMIAZTJAncNjsW+GvNDxsoNyYWxgV6ziO7iZgKba6fNv2GtCnjQKlcexrGx83NcLRj3AFSJG3gfh6yrPLuSWHcdq0smBLcco4VrhEKm7gzVkeDqxdRVJM2xq0pBHNiEhXdjACKdhQZ1HghgYJxVzCxUBaBUm6BcEf6TTqnMzuCu3L9NHBz8GxkyuPh5mt8VquxJgjSlnUUSo/vR9aZBJ0hIeycjTkFy8cqxk38asgbLbh9CaAbQoi6cY2yy3ptPiTFvCoiZATsISPxsEx86dq8MNxqtDwUijS2sidIQx6GhPb7hCkNh+OIJ1fAEa6kpe3WFgz6XQMxNHHz7kVFChh5aJf5aLgjIk258VOVfvVkrbj8k5HttDdwNzK/0uEEL7qG6+MdvFyPHhtZTYk72bgNIWI9Sr2xrMnAuN7SwC3WSatf5U7S63J60WgVw2rpU7sZB7fL1GGOI5LcYnL5ujZDcbOM/xFulnchE8ncKBlw9qxqSXap2IJ953bVdQchXoxe0+OKMmtKaXR2hL6J4KBet4gCXCgTIKHMbigSsrcvjV/5RkwKRptGt+z9LVLRSsxsvJKlGP2U7rs6TWjiVmIYM3tsKbZmLEKDm4Il+h1u4lsCq5GTFw7xtK9fmcmrFItsh3EnCyLcQLMoKREJaGSjgdcn2HFzrBl3CICuECRaxvHpDne+3i/tFtw1/fa4uS/JhsviNhfD23Dbqt6i5tSaoYoTpgCp/A/uXqHFYyTcAOk5TZU7efOKzGpc3LrrGeN2dHJGpmmQttVNvClmJSSNlJkJWpugC3gykX43pQir0osyZrRcj4i+j9TOGMmAjEq8pqa2xPzcNrk7FYBhkQzFBCn3+U1xmrjdE4qa3sYW3ACPf0unI82roVP1Ota1+VgeJ3KmEALUGIgWS2GD8YiyOoS0UY1rN9iqyNSURKZMZ54ClEfcQ7m2JiuszWRlIwIK42uZMaHCnfJDGZwN3uGW8TfjrsfBna/NeGNNmNQIrLgXi82Dk2jGLNfS2o7wzK/PGR938P1pwRDQqV7y8abbxKsSd6AAzP2TvOt6DCEE1HXtdU5/xYzbF/zViRQ5ZmDakHjTjbFG4E0/5CLkIo3+LSPK7G1cWsT3C4uL1I7TL+rDgXZDmHyNGLmribQwXNquC6Mq6h7MpManwC1M33betth6i2nWhwrYmIkQsG71aix57BmEEPCe974Tj91zC37xu1uo7SZuv84E8Kl0C+3Kl8IhIuBFhx6G151+BD72kU9j5QBjQgP39Jmz8ILttqL2zelt3jyExx5bhvWbBps8EtxFcDFqAjlTui7kPkKwInPowfs/eC4euOXPuOza21pwx+JbTpEhugAAT1eZltM1Eyf2A3EMA4NDytOyThW4xqWdR/oZKQgJKzKfA+mK4i6Ogc6h4KnQ78wr466LwAmoHgWHm2214I0GCFnaYPSEyO1LqwFdSVuS4xtzzAlVV2n2jA80Jy7nskPRLIG8Y1EQbGx8QgUuyHgqUJ8abVhwufoPuGjNswXplI3RmitGeYhhxxPuqLhPfNkpOPuUg5+3jgEAN1/7e/znZ38EIGD/A1+ICesfJwzwuIkGccjNaT/GLQpGuF3UDZg5awvsu3BX9PV0AYyqUvqH1tK1C1+0Pz7z3rNQuyXI+WwIGBrYhJ9fchkuvPj3GBnj7CL32xIg5N7GI/sB0M1rIhRjCF0ceNB+GF3+MPy6kTx1r9PhlG0oHyogyGZLunhfHXCajWg6W3Fin7zg4+hbsxTnfvRbzelrub6t/sGpCAU61XvNc6UOSGsddOgquimyjPbP4WZjFRoYt+8nqUOR0SEkx1UOrXSFsvRNDqzNaSEgTZ2Kk+AIrcwoeAhAinjNBgVf2Q7FnVBkHaRYtjs4W1T5W6K6pJEZHBV53FieFKSxfDmKcySGuTUO5K2H1+GMsz+EUaf8lF2EgJHhYUXyi0suw4qHHyTcVWFEhql4FhPNzzi4EfIwxjKixPKc7kpK3sjyjA/vf+9H8MBT61zf/ZMm47gXL8LZr30VZkzpw2e+dannG8u3yALKPS5sDQvfI3eM4uKfXoYnHljiz2kMIjlyNgd5IEqcryxoyzQI7rJw6dbPWKDTPUXLehEXORvZjsdjhs/OPF1XLiz0AYN1j3Dq7WyDFsBkmt0KlPl4W7GV+NY47uqAck3TcQbE9CqA5KmKtsr02H0kMvgn2poE0hSdgOQiKWDXxPw0nEQJcToB8CknOaEcxYJTZKYlGuNDyQCZC2fSiXHkXWOObqtXr8MI8E/gDvj5xZe6cbtmMCFAVpeWD3k5g/xncAd6uK78uLoN4Yredaxfuw6rVq/1965eh+9954fYODSG8846Fddc+1fcsXQ59AlH16ZlTo53UpsYD3cAEMdw8c9+Tc4k5Fs52+MIDpV3E3cZnEKBm+tTPso2l2NTRlRmwq24M60ZowWsJm7NesBZJmcmua3osznV8wCoM2JHof0B/slXdngtTrsYpnodJL4D6Kp5ciGsbeqt4Z2aHtOBdAxlQouPRvIcHVQwRYbD7RFtrpAW5SGgAL8gS241Zslc9z+DW/WtxM2RJ/cte1nMnbs1hgc2YtXaDQACeib0YustZ2LF8hUYHkmPes/dZi4WbLc1KozhvsVLsGrtplbcVVVh2223xpZbTMfw0BAeefRJbBwchhbGBLcoTKyh772I1p7W6GmoEB0OKH8QI3596VU4+xXH4sXHHIg7ll6O0Olg3tZzsPLZ5zCQkijMmDENHYxi5ZqNyt8AYMGO22PeNnMwOjyEh5Y+hmdXr4czojoCoYOttp6DoY0bsWb9xkymBZlOt4sXvGB7zJ0zE8NDg3jwwUewat0m2NO6vAAtfXp6JmDnnRZgy9nTMTw4iCVLH8VzqzdkXxbQP7Efc2ZNR/+ELnr7+7HdvLkAIlatWoONA4MmaBcsKCOUTDTawiu7sAiExmDY80IAUFFiLk6QgitKeYiex3FxE7H5awxaZczZV3N6OcJtmKzD/6aDDWkYksOru7ggumHn7HUKI2PmOSfGBHIEAv2O8EZOBqDt+chqwBKzg4x3G4Up6VvwieMRZnncFgFtFZ5MtzrPTFiCZFxVB1/838/gnt9fhvO/eRkAYKsFO+MnX/kPnPP6d2DDhNk479xX44CFOyKEgKoCBjZswMc/8QXceOdSxd3T24eTTzkeZ566CDOn9GLV6vWYOn0aeqsal/7qCnz7ot9idCyv6nR8lcfLqa5U1EMCj5+LYpng2bxpDZ5eNYBt5m4JAJgyZ1v85ML/xoff9xHct3wE737H63Dwvjvj95dfhvO/cRlCAHZbuBfe/bZXY5cdtsbo5hFU3S7i2Chu/NNN+PK3LsbKdZtgUbuDr3/jAvz5sovx+e/9luQAHHb0UXjbG07HnGn9eObZVejvn4SZ0/px3R+ux1e+fQnWDWwmmSTMJ5z0Yrz51adgy1lTMDy8GRMmTMDY6GZc94c/4kvfuhjrB0bxwkMOx2f/8zUZ5Bb4yYX7AQA++4nP4Nc33Jf4oBG7DG4+8wvlCtC2TCfkl/RwfcINddlYi2ClmUHuU52YX75mmVDIJhsgpYUQa3uOxGVAyVnbCIACX5ttB8SuUhdp67hyiODsIwNw9lIUp9iAG0tqswK31AbSLVHbUmFwKqnFMe6TaHUP3fBHaC5SM64D6CcXfIvxYyzHcy7TousaGZcV2xbstgf+7a1n449X/x6v+eLX8Mxz67DzHrvj4x96G97776/DrW/4MIZGU1vHnPgSnHb0nvjm1/4Pf7njAWweGUWn24Ojj1uED7zjXzEh1PjSD68WBhgNSpLIih1G4TiF/+y08+nQ7ceMqb14aL1lDQAwY85cfPW9Z2HZksX41AVfxf0PPAIgYv/DjsCnP/BGPLz473j7O76GxQ8/hZ7eiTjs8ANx7pvOxDd23h5vf8+nsWLdoAUmJUeytYDTX/VKvPM1x+OiH16Mn11+PTYMDCOEgJ132w3ve9eb8NUL5uHt//k/WDcwonS97pw34E2nH4Grr/odfnDJNXj62bXonzQRxx53NN76+tOw3TZz8Lb3fwl/ue4POOpP1+GzX/w0+tY+gnf+9/8BAMbGyqyA5crHCnmrsQVvJ+IEYs2aYZE/76wWuI+GThe0qDHLoSJjlyymLpyPq+EFu1dlX2BUOzGaYow5s5AxE4o6BI//AlLKLpXaFqalbcnLKZfCGMuZDclqNIWNmd4WwTR+F8wt6El952khdUrllBO9oo/rEMTAlHR0sOvOCzDayCqSQ3x62TKs3zRUkFg6wYC3v/Us/O+Xvoorb/y74v77XXfjOz+9Gh/8t1Oxxw6zcfuSFQACrr3ySlx7xWUYHTN+jo2O4A+/vRrzt5+Ps04/GT/+5XVYuWmz74+VxBXpCqVx3xRJ8rF9DtgPW03txY9vv4fuB1579pn4xU9+hJ9c+VcdMk6eMQcffvfZWHrPHTjvI1/F0Egaf4+MbsQ1v/sDFj/4OL71xQ/gvW/7F7zv0z9M+4kV9aGIiO133RNvf+2J+P43vonv//rPSnuMEQ8uvh/nvfd8/N/XP4m3v/YknP/NSwEAe+x3AF5/+pH42Q9+gK/99FqV44b163HpLy/HUytW48SDd8bMaZPwzOpNGB0ZzfGqxsiIrBKNDmMjS2gM1eDPl04mij6LLtNT2eDXVozzccMS6ZPbhv/NGUrwQZYXxjnHpZlDlYfjLbjVLhG6qCNQ2eIpXoraTIlgT3tGP26Sgo17KK0cWpSKK3/XTQfiH3SiaC1j75AMkMwRzU85ZADKlM92qs4ciOWUW0Y5YSq+9uX/aukjfT7+4f/GtbelCGuOPmOnqH3LDdfjyhvuaWQtd95zPxBOw7bbbIXblzwHBGB0ZLMWtpSuTPPNt9yFN552OHaaPwsrFz/tnSsVGH2BL0DfH8voouzgbEOTnXffHR867yw8uWQxfnfTffmapDgP33sXLrri5kxLouslJx2HGX0R7/ny9zE0MmayyfJ+6tEl+N7Pr8V5Zy3Cjhf+CkuWr4dzWFnmZ5x+ItY/8yh++ps/Q+owUqyLiNi4ZiW+c9FV+PA5L8G3f/wbPLthGGecfgLWPfM4vnOJOAqOtjVuvfFG3HrjDc3InbFrMCyyQzZ0IPLzb009Uf7K9YXeBsCCUW5P7aTSNrxNxYwbNuwIFkx9YZ8dCGGKeQFaq31QAC8yvJYHNWIXVSheAEOZBGBZARcBc3oSXGFEGCD3ScokbbKnjPpfc2ZcKMrXBsCq3+X8MWwxmeKKXogSWbldbT9QFmVCt2Bn50IIwNBanH7WBzHisutBU10AACAASURBVA67d3BgQHE05vfp75tuvoNoMNzr1m1AjMDE/j7DHSp0Oj3YYcftsesL5mNSfy8GNm3Ck089g6GcavZPnFjIQLC2T9O6yAPgY5/8MIZHaodlwoRebDVnJh558AF86OP/i+GxJA9p/uZb7rColf+737574vEHH8DS5euJj9JP0pk/3fBXvP21J+CFe+2EJcvvUNqU6s4E7LvwBVh8x43o9k/CZFevMoVfvHgJOv1nYuHO8/DHe57G3rvOx23XXYWhEV/vMoMy3StH+zystVma/Ch/6NjV6oc9blXg4PVBZdDI8EgO0j8Vx4PWNSxjUKerx6LujQlkxyWgpPAq9OlIgPhQrrnQ09xnM4tJq67K5d78SgAaSzqQxDL70whx+0m4aRxzTKHBYDLizOxxpwYLIEqCu56zm6ZAG8vcqV1bFmup4/r1GzCiqRulcA531cIjiwK1rjCtkQpMeQ0ITyJlHNvusCM+8O43YO60Cbjljvuwcs0GzJk9C0cccQh22nG+YQQw7tODlMlpTSq/6xIA7rz9Ljy3bkivQQgYHRnBIw8/hpv/djc26xCIom7tA0oIATNnTMVzDz+UWd22YA9Yv24dhkeBmTOmufaExm63iykT+3D4ccfjymOObcqFPvXoGKZNm4Kevj5M7O3BmrUbqC1JnQNEzzSDbB1C0JR+5GhPQUGK6jRtKZscRVeno3Zd0d/rYiBDT6wsA4wiBSTL5g/pOS9JD5KVIwe8Usf17zLj9kGfSUEOwN1MeT7PyiU36x3UMKW47DFlSksYq9M9xMUoym1KbLtCKfR27ydMivy7qZQWBng+mo7L78ZUUnG/GrocjZ6hlD463LCdwZr0d8gZslC4T6Bv8gx8/vz/wNLb/4z3fOWnGBqtSUYVFuy5D370hXdDZeWGIeKMAJYdv89D+v71pVfg70+sNxwql1y912hL/GG55ki2fsMmzJw2NblWH7pzlxUmT52G3i6wfsMmz5N8w9joKDYMDGHp327BJ772i3yfPU8USK9ijBgcHMRI7MGm4RHMmjkNnDFR40X6T3ynYq7pQDGNSGCsqB6Rnixm3gj/fUDyu1h5A21/tw3RJjyXwMQYEKEycjNbcq0Eas50KGhqtlPOfDYDcKppxPzCSwARNmZN97LiFOkVex/+rZeJcrZ0nE/reN4aTSfcm6xZ+XPjDcdj/WsEYYNuLUyZg/FjP76+iTs0tjeLpmiKO6D5cl5VF6Sxf7k5avQ7P8eI3ffZG9tu0YcP/uDSIr1ObYyOjtm9oiDR7vePLRffbAAcFFxWJo5WvgtHW9B/998fxJteuj+2mTkJT63eBJZLIqnGwQe/EF2M4e77lrpmtGI2Ooy77nsER+6yIzYPbMTASFnNbxojMIK7738cB+y/Lyb2/BIDm0l/XMrtcbu/G4XEQG2QrpVDCf0q7IPON2WdEYu82jLbsl3GwAYdiT69VoJgEdwVD+jZnObS8EZmoYkBUNnDtOZtWvelJGW3oUluLJaXsdLxtwBvM2DussUDR+6EQBCTGtu9cz3CXQ+9Z3zcJX6KBKI4zjgFC0ei0qsLbW0KEvJlWcnqFDWmTOknuk3B991rVyNP+hd9UMNvYij7jkW71Gj+WdO5gv8UsX971bUYCn145zlnoMvPJ+RrZs+djzeceTwW33E7Fj++Cs7J0+9f/eoqTN5yHl596uFFP+lfp6cX7/r3N+PgvRdoF7/41e8wZct5eOO/HItG0TECC3bdA5/6yLnYZbs5jgW2oU6hW3ovFeaZY/on6zAt0FKaA8mbrlV5hdxeLPiZeS1Ov6TLZR9yX5PnTtaiVw5TKdeIRtDJ3zGmeZAUFhtj7aIzbrT0rsp9uU5SYB5iEPDWdIc8tyuO5qZccVRSKQLdRnug68g5RXZYramrj16KspFRUT9yJWGzDWLbnBw5MfL8kkouvvsePLNmCG9/62sxc0qf9tU3cRLOfNUrcPpRe2BgJKb0O/c7NDSMGAIWHX0Ipk+biq3nzPQcJtxuU1/HP6ZNF+SgaKjhjFYuexz/8+1f4aCjj8X5H3gjtp87C4gRnZ4eHHTowfjfz70PvSPr8Zmv/Di/hqmUf5L5I/ffi2/+5Bqc9Yaz8cYzj0XfhC7kNXyz5myJj370XTjuoN2wfMVKbWPxHbfhuz//I858zavx/re9ElvNmgoA6O3rx9HHHYP/+cQ7sMv2W+O51etz1AUGB4ex4667Yu9dt8Ps2Vtg0VEHoKMiqU13lDyTN3NOvyXYlIG2Tc+LABqk/ZLP2ek22yWeKZ3cLsjRBIfFFrGVNpz1taSDglu3ASLQo+gKiEFyCCt4YHvpkE0FS4vckEUKfSiiLrwzUe+Zx6pZ0WytfEFEsVLRHJXBaUw5aaW8xB31l9HClwid5GjdOFA6LBxKybhgb5MSzz+8aR0+cv7X8ckPvAU/++EX8eCSx9GZ0Ifttt0St/7lL3j3Bz6Pr3z9c3jlGSfi579PMyx33noHnnrupXjz296C179lDI8tvgtnv+eLqozkejWD0ZmmjC3wMErSeFdRZzn5BXfXXH4FBjduwL+fcyZ+eOFhWL9+A7oTejF5Yi/uvfNufODL38ejz6yBpti8NQKNry/+0UVYt3o1zn3dmTj9jFPx8GPL0Ns/CTst2BZLFt+Hd7znfDy6fB3pSMSPvvsDrF29CuecdTJOOOnFWLdhI/r7J6K/twe33fI3fO4rP8TqjZuV/ssuvwYHffCN+OpXPok6RmxatwaL77oHz6wdyhlCrgcobNL9tqxNgy0Fg3IRXDnsCR63qUbQ6+0RgjLgwNFhbxqjcoIpbhNHowgtwbC8Xn4GhIOPfvlA6PT1KxFuvCfUc7GRI6EZlDfe8tqisuwcgU3F+gVbpUf2H9uYxja2Dc4pUV+FIUuFOJROSXHL7Unwc7baCrOn9WHxA4/aFv6KQ/B5Bdpp5x0xsG4Nlq1YDSBgQl8fdtphGzz5xJNp8ZY6r4Q7dCdg9523w4pnlmPl2o3a0oS+frxo3z0wZ9Y0rFuzBvfe92B+DgOYs/XWmDd7Em6/92Hlb/+kydh7jxdgdPMQlj78ONZuGCTco+oYpkybjvlbz8KjjzyGgc11ZgE/l9OM/N0Jvdhlx23xzLJlWL1uUytuxIhubx8W7rEz5s2djZGhQTy05BE88sRyyo7lnh5cevl38OfLLsHnL7wSrE+Cfa89d8E2W+ZnQx5YiseWPYdaZN+yTL23rx97LdwVc+fMwNDgAB54YCkeX/YsnJFnndhizhzssmAeNqxfiweXPIHhkVHrX3Rft9yPpnOMW/SkqI01N8GG79/RP84nylomW9ylNubsyt8j5931fK51GJwwuuxecUdgbHgwHHzkyzehO2GiG28FiT4+9ZHY5MVTpk+cfRROgXE57zyeYQsw8fKx5dpICp7+Njrz032FI7GoihYB8gNyuT2ZlpLcw2UYbRnDeLhLXsnlkYTDNHGW5A3J45bbUhuG29PqntBt4LZso9mekM30F1gdfSIzIb1dOadvtR0u/cEn8cOvfxPf+/Wf7V7OOl2GKEYwHu5CLxFVnv8s7nKQMT5uf4X9zouaYnq/qn8hc6nj8O3qVHymzwWtdI2uNoYt6rL1oMFoVT1QJhnuQHyMMd/yD2y73jzYtauaaY5Lf9gjsRLHCJlGSjSmNMjmtgMBL7OWIh3itJZkImsInHGQ19bpqcgb3ETInHh6B1FeaKMwTfn8R+4jmmRhjLbP99uKN8PNfCSGk7dGg7eCOWrboepIgkjLcaEC1xoKKUAabqTfQWlIMjKEseXxmZZMK6fjgduPQigt+mIFV6VnTOl31e3BK884EQ8uvh+hdyLe9IZ/xejGNfjtn+5QmSWWd0yRJSsS+Qm+VtxQ+pM+Cj3yNQ5uJTQabspc0wwWlN+2OrVwaK72JOeKmlirjufFjKGJ2yYEqiyjKushr3YmEiAvM670BUfMF6YzxGgLMjPuUNN2ia7YKY+oa1rFDcKY55DRwy/ZK6liqiDLe0DjXqjRJT2OxbXsWKJiS8eLSOvGiCLMhiSgK9Jyu0G8ajGUsuvZv5YOJTocYNyuPf62W5u4UfTPuElSDhrN9zuo1L8bigluIbcqzlH/YTzcfJhWCOaUVfdnkAIZZ0q53SkzZuGwww7EW84+DVUV8NRjj+F9H/wKlq8dBPPb486O3/GWl2jDY82/AzvITE+jVtUY+4uRiIM1GgINNUTXEeBfm1LUMvyqUMAFyYZqML8Nd/qWwNxWcDZnqbjpVGOvjsLBpuuK2qHQ6NBEhIOPPmMgdHr7Lb2DRRj2MBohxLNSup4jrz3fL1He7+2njMhK5dc4oLhO/oYdaxunubGiATYsRTuR6UzXyx1tS8odc/WQrVJ197YqnyxuqlvOlU6lzXGKYyz4Mw5ugLeUs3bF4ZpMZKo5eB7pLYbbNmvJjz2DSsEuG2kZMhU8CaHCzJnTMaEb8Oxzq5Ee9hwH93iK7g5FpyWhMASrpeWiJdupw81GZEuw+ZzT1SDPxQB+iEzZ9DjDL8P6/4+7HDYHWQ3cqFeY7rkYrPyJnmeRnw9Lq4wDgFgPD+pTp8l70lidCjtupWKwZwTMuCRNs9QrhJIRME+bGRqyosaaN44pDM49fzLOIpJYA1VHZa8vZWnUH1IocPsQBKSoAfLg7Palfeo7ED9Sn7yAqWn4yakUxbgAxFpSZdj1jtdEA+iyEBxdso19EldZPRcjLZ1yADBGETs3zsOHzHML4Db0tF2bGHcRLvma/CMiYuXKlUWQQHoZjltQZ/cYb4RWcXK8+JiVXgHA3rMbIbN1QbdTJLrdDII4h3ysCgVtkfjh8ZmeFTyIQIxjJhtJSWQYoEOBQh4Fbp7psJ3WOv66ANLxiPTu3JyZoEO0+fakDVvSngKLBJVcDKhNOdVIjWl2QFDLvG/6Lc/mK2j+kLHqugNqM4oX1FmI4PuUlLnNUcDaS7qdgQV6vgTpt0Rae3cI0avTXlbQtchMXjbWsO3c7a3wz/c+VWgGxnwRPrFxFlNvzgHRfaHAnSOcOchsACH/1ohOETTfb2+4Mtoaa0l0xWlUuu1JXVpZqBH6+Wa0aqCmWTP9V86EwTst/ptoi7HWnm0s7x86bMNtsxktS6jVd0fDnWUvqy6be4rmAEhOyn3y/UE9uhg1zTg2ZpboOqU/IxDcgdbLhECO0dezzKmUReOCpyVuZ+sy020hmW7Ov2tSdPY+6iGFCIsczsBU4ag6rmBSnzrXX1ERR428ZWjgvLhgjOjr78Pk/gmmGNlxRFVwoH/KNOw0f47hDAH2smej3c0EkWJz1BaHFBzvpF1hPE87N3EjVAhVB7vtvgt6u4xbFCqg6nQwe/YszJo+hfM0xc08sKJUoGgi1xldJAwypAJ3xq7yjRFVtwczpk0hqNSWjs/rtGxflV1wsyOoMHPmTJN9gduyt4xVghcCqk4P9tp9gdIkj9kDwLztt8OMyRMARMyaOd0HKDcml/b4Hzu+gFmzZua4EommNt7lP2sxrBK3GTSqSh2DODZ9pgMYR9+FZ0FpUedRDo9zyUBXhWrqJbRSoGoEMWS6OsXfFVDHmMYLOQKFyjyTfrdGOHKQORsIbEwcOVyLUZsWIYaqA1QdAxprZYAZeeGAWMAk+Fe99tV4z5tfBmjqFLPS1uphZ2+7HV56zIssoiEAoQW3E5JFzhgJeyBlUP6U0UG5le+vHW7EiFiP4RX/chom99g1Yuj7vOhF+Nwn3o2zX3kSzn3r2bjgv87FFlP7YRlb9O2DcEvqLM5NFo9lp5y+i+zmeTBEREzdaj7e9YaToelqaQxZ9hQHm7gRMGHiFHzrG+dj3x1nuwxNcMcWhZa6S6enD6975UsMt46zI3bbcw9sOb0fCBU++r5zDI/IW+VOWUTGbUabePLB970VEzrywFgRMADKUqWd8XBDcSd5jOVz0XTc6X6JW9rzxu1XR4+ZTnANiWkuh02Mgw679gV3FUI3jo3le/jpvMLbaJrILY1TmZWPbmhDwnGfZICNh80aNQJhVC5QGRJqBZgwcRrmT60xEGZj1qQerNo0YrQDmDS5H4MDg2o8sR4b34sDmNDbh24FDAwOg1+iC0T09fcDY6N5EQ/U2CZNmoiR4WEMj4xShEybxNYjmzE8KuPeNIbs6elBTwcYGNrs038kHszfeXe89pQD8JH//gI2DacFQzvtsRdOPvZAfP+Xf8zwKkye2I+NGzd5DueMZGJvDzYODAGIqLod9HYrDAzl7ehkLNrpYmJfDzZuyo+qB6DxqocoT3sWssqfyZMnYmDTQH6PDi8nl2wjHRfFP/Sow3Dxjy7BCScciTvyE6aCW9vNkbGqKkya2IcNGzZCDT9fP6F3AqpYY2hzkvfVV1wJgLddzATnF/NM7O/HyOYhjIyKk0zEdbpdTOzrxYaN8nYmKA1aXynqZvLMUoqXnEkAVaeDSf29WS40BE9CI5weq8pFM6FY9D2OjQpfOIjocKl4wJJrYRFkg17mbjiHELsaXcqOmSjnRIigRpWWCHQChzLSvGGgbpjYkikMooLN/2WvmK879MjDcNMf/4Rl9RY4edH++MHlfwEATJ21BT78H2/CpjWrMIaAxUufBkKNOfN3xltO3Ref/OrPkSJeDz72oXNxwee/g7PPPgMYGUK3tx+TwhA+9/VLMG2bBXjjiXtjoGcapk/swY4LtsP/fvFruPOhpzFzy63w7nNfhaEN6zBl+kw8dNet+O4v/oiJU6fjHee8EsMb16Pq7cPAqmfwfz/5HeoInHDqKTjp0N3w5DOrsGntSvRokBJ8Aa94+Qm48Ls/yo4ioV1y39+xdHH6vd/Bh+DVpxyKZ1euwZwtpuHC71yEvz+yAme/+Q1Y8/hi7L3vXpg0dQbWPvEg/nDPcpxw+F6YveVWuPPG6/D9y27EWW98A8ZWPYGddtkJqHowZcIYPvOFC7FqE/A/n/w3/MeHvpTFE3HBp/8TH/7Q5/GaV56MXXefg/POGcNXv/1LzNtpF7z+zOOwfPmzmDV7C9x64w24+s/34dBjj8P2U0axYLc9cesNf8TVf06b4aaaUgdHvnAHfOrTX8e//8fbMGtSF6s2bgZCB5/82L/jxr89gKNetADnf/bb2P/IRTjlyIVYsWo95m45E1//2oV45NlhhKqDV531CizYejq2224eLvreD3H97Uvwr69/LZbc9DvMXXgwtpu/Ld533uvw/e9djKHuZLz9za/AxrVrMGHiJKxZ9jguvOT3iCHgpJedgqNfuAAr1w5gy1mT8eWvXIgFe+2HBfO3xrve+Xpc/LNfYft9D8OkDY/hNzctBhCxyz7748idJuPbP78Bn/qvc3HznY/isIVz8bELvovDjz8eh+45DytWr8dWs2fgRz+8BA8vW+V1uaUGo+f1Z3ZAYkdqZnVhd2wqVPvidRquD2rH3QsN8uVCRoQQuq4AJNNLkqLwTIKMfWQNAnu/YLMO9gRh0EwvZA8Z5dl7HucpodI+FX00byiyGrlZrqu6OHzf7fGZC67C5vpxvOal56Jz+c0YQ8Bb3vJaXPrji/CX+54AEPDqN5wN1M/iuacewYQ5p2F6X4W1QxHb7boHnllyHwaGhvHd7/4Em/Mekq998xux/25z8dCGCocedgDe+Z7z8cRzG7Bgz33xqkUH4o4Hf4Xz3nY2LvrOd3D/EysBBBxzzCGYUAHnnPNqXPXLi3HvoyuBEHDsSSfh1KP2wt+eGMaL99sW73r/ZzESgS222hZf/ezRkMGCfLbdYjIeXraaeJE+dV1j+pxtcPYpB+D9H/sCBoZHMXnGFrjgI2/Ge9//WVSdDnadvwU+ecG3gNDBV776Kez81K/xyc9+G93eSfjaBe/Ejy67IUW/njF84rPfQozAwv0PxHlvfjk++qVfotul3cFDRKeThoo/+tkVmP2K/fGlb/4c3b5JeNvrT8bHP/5lbBgaAUIH737PuXjwoUdRhYAD990VH/zUN7BxyO9zueMeC/HUg3/H5rGI31x7G0465kX44RV/BULA1NlbIay/Fh/4xDXYZsddceIB8/G+j3wBo3XEjDlbY5e504FnV2DbBTviwu/+FD95ZAVmbbMDPvKm43H97UvQqToIAbji0iuw6ICd8Nkv/wBAwPs/+G/4+fd/gCXLVgEh4JQzzsBxB+6ChzdNwkELJuN9H/0S6ghsNW8+5s6chuuuuRYnHrM/vvCV72HzGLBgv5BfXJZqMaEK6FRJLltssx0Gf/t7fODXV2D+rgtx8Aum4uOf+z/ECEycOh0fPu9f8V/nfwMjdbSEgWsJzhgiswriYLlGaJZNtqgZnGUTrgMO7OVsmUtqU3t+xXMNxLHQTVtyifeApZ9S+UW0Ybt0So0KIF9pFWL5xSjZ6Gv49EuBcNZgsxvJmXWgU65uejVlIDvusRBbTevDKSen3ZU6/dNx6N7b4abFK7DDzB58/r7HIRnRTX+5E2ccuA0Qa/zmutvxkqP2w0+vvh0nHnsgrvjxRQgBOPKYIzB/zjRsHhnFgm1mYtWMqcD6zbjn9jvwxLPrgRCw4ukVmDh1IfqmzsLUuB73P/GcCui6a29C6EzAPrvOw5ML98FOC9NMRc/ELvbZcx+Mzh7EH66+HiM5NV65fBnuf3QF7AGmNOU3PFKjf0IHgyObbWox83qf/fbBn6+/IT3XESpsXLsKtz+8BnvsMBsAcN2fbslZwRiWL38ON/zlTgARo8MbsWEwoqfbQUDAHXffr7WAe2/9G17/L4vQ3yEdQDCRqpICoaqwzY47YVpPwPHHH52UGkA9VuOg/XbDsjrgphv/io2DmxuZ4stOWYTBZUtxxsuOA0IPjjlmH/zkN3/FaIzYPLgB1998HwBgv/0W4rprb8JofkfommeX468ravRMnIZljyzFvY88CwBY/exzqPomwn1IvXr6J2O37Wdj4YteiL32T3j6+irsdODe2GLjRPz2t9egrpMNLH/yCSz3gJUFXK/gPgbWrcSNtz4AhICDDtgXo2MjOP2URaqrk2bOwbxZk/DIc/QahEivmwDgX+BUO57pEFXsqKijNYxdP7GwFTpGQxx9QLOlJKCOClXsupORes4G7Nc+II/9QnGP+5F/y9815Cl43jXcFsrAHA95Vyv68nHOaKy3U088AhdfchWWrUnjzYeeWIPXnLQIN913EWKni55OJ20PF4CqqvTW2266Gad/6I247OZHMKszgCdXb8Jhxx6PLaq1uPDH1yPGiJec1mM7SQp2KhqOjmxGt7cPFQJqrkzXoxgcGMRtt9+DUTp+7TXD2PfwozFj8kTDA6BSD16rN//T3+7HiUe/ED++8hY13BAq7LbzdhgaGkb/tIlUGwiYPLEfQ8MjwmKIMsU6JtqNu/qr27Xdz6ueHvRUwFhdI+R1K6mZDvp6J4CVKcaI4cEhrF+3Frfcdo8ev+W2e7Bh3XrsdehRqGX7PllfgIDJM7fE3L5hfOOmu9QoZm87D4csnIcb7llmRU4AA4NDmDllkuIQXQkIqGte1ZmwaMGRU3oA9dgoBgcGcNvt96aaSpbh1YMDOOzFJ2LK1Cl5vUOuy+jmMAoWsY7o5uwqhAp9vb2q5jHGfE8HmwYH8dS6p/HX25Zmcivccvu9eHbNoPJNDN2G5BX9RjNwk/5bLUZ2lBM79W0zv8weqb0AyLoT3fpStnyk2okMgWKsUTlDVMIoJSqnV3SaNFjDXDBRsPKv0lmWEDr6LzWf1y04hwDfltDG/VKKNnnWVth20ghuvOMBLH3kcSx95Ance+ft2Ng7G9tM6+KGOx/H615+FHo66R2eJy46CJ1uF4hAPTqEux9fj3PPfin+dN1NQIzo7etFPTaGGGtM6OvDXrsvQLcrr1cR3B2lb2xwA+5+YgNefvyL0OlUmDR1Gt513usxZUKFP9zyEA7Za3s888xzeGbFahx82CHoDaO4+cabcdQJL8Z2W05DCAF77LMPdp4/C52Or1hfc+Vv8YL9D8fLjjsQkyf1Y8asmXjzv70eh++zA+667Xa88PAjsMPcmQAidl24F3acNor7n1yrMvRTaX4oJ4Z2ysnHY/qkXlSdDk4+7RQ8ft/d2Dy2GZvqXuy4zUxUnQ5efPIJmDOlB91uMpapU6dg8uRJ2LDiSayrpmFGf4Wnnl6BlWs34aTjD8PA4AhkSBnyNoLIsxzHHn8krrv6D1j6yBNY+uhTWProk/j5pdfgpJMWmQ7kCP7Xm/6Kw447DvPmTEOoKuz5wv3wmpcdAQloUdc+WBBK6U1yOL39/ZgysRcTeyJuuudJ7POCLfH0M8/hmRWrcMRRhwGjw7j+uhtx8mmnYMsZExGqCi865BCcfvwBAIBuTy9mTJ2MqVMn46mnV+CF++6BTlVh5uwtccpxB6HT6agehqqDEAJuvP7P2PeAA7Bp/Xose/pZxJ6JOGTvHbF5dIxsiZ0ZZ12s53QJ2UNE3Ypbj+WrfD1C2iU+6XU0lGmbLdEyBWJn3g57fCh0enpCmS00HACnX2zI8Oe19tCSDpW3STXWjdZlkZYQGRH1YSYBmh8XDgG7L9wdjz+4GI8+vTp5wrxhyKr1Q9h+zkRcefWN2H73vfDql78Ye++2Pa666lpsPXdL3H7PgwihwpPPrMZR+y3ARZdejxrAk48/iUOOPgpHH7IPdl4wF9ffdBu23mIqHnx8JWZPmYB7H3wCQESnOwFbzZqEuxc/hrvvvAe773cA/uXUY3HoAQvxx2uuxSNPr8ED992P7XffC6eecBgO2n8hHn/gPtz10JPYPDiAex5ahrNf83IsOnw/xE2rcONdj6LavAHPrt6oka8e24ybbr4dO++xEKeffBT23eMFuPWmG/DrP9yGkeEB3Ln4MfzrK0/FS449BPNmTcSXv/kzbBrajNlz5mD5k09gzcZhIARsPXcrLHngIQyOJt7Nn7cN7rpnMfbcdx/cdctfseglJ+ClLzkS81Fy5QAAIABJREFU2Pgcvn3R7zBa13hs2Sq86XWvwIH77YFHF9+D+5Ztwuj6Z7F8+SrM33VPLDpkLzy65CH8/k934MSTj8cxh++H/ffZBdf+/gY8u2Y9pkybhrGBtXhi+RpTyNDBEQcvxOVX/QkjtTzyHTGwbg3m77Ibli6+H1tuPQd33nkf6hixeXAT7n7wKZz1qtNwwjEHY+70Hlzy62sxPBqx7dYzccc9D6VMIFSYv80s3HbXA9hizmw8t+xJrFo/iNg7BWecciQ2rFqJ3/3hJuy5/4E46diDcND+e+GBu+/A/Y+uwNDG9bj/8VU4+6zT8OKjD8KM3hq/uvIGbB6rMTjWwZkvW4SxgXW47fb7sMOe++CMk47AdltPx09//jvsuMNc3P73hzF/3la44677UceI4YGNuP+x53DWK0/BIQfsjR23mYHLrvoThjaPql5bfS8HySBPxoo9sxOgBwJdwtAc9vv4WtFxrlGwbVJmFloclHPe9Wh+NiTvZ9EYDgRw/cDOy6eGWzLrnERAOfbysyfBvB8VSq1vquS6TAQt9xRtKeJI3/wpx3wBTU9c4BZ8NEQzzwzP7BhTjSE/weffMcG05hpFDHAPrxU1GX+soL3Rf+GkwZf7e88+501YfP3luPWhFXqv7Tpd1IdKHtIslz9mRfLyKWB3jS7YM53Q5zgq6rdRI3sefWqj033GkTfNOrgHv1rbK9J8h1uGF2Mpew5w79nxU6YtMqw6fhFkibvBsxZZ/9O4Qz4UWjAD3raBODY8WEk0T1+8qEM8Um1Cj7I1f4S9PEdA0wIdrc4yBTTGUgyUjZQr9tw1EYj50Vk3e+NcbcEYboeGENoJK7AU8sbBLUuUeUwpbfBiF0mDRShMQxtuwJTKCYodVOEMXLU7eJ4EUwCHOzBu7kVSUIC3FbBps3LOHtZuyDJnbKURONxCi/xsrnEJ0kZk3NROmdG24hZdKo3JUJeOIrADz5c0cUt7nJq3OHXWLXbSIdMnmXe5jiWEvIAwEm+8M20OzWHtNnQ8NHWKMPKrOpyZ6rWMJa82PeToMwbQ6e03hkS0e+zi4+Z6+T7v+UPFVd7iPAN3/ZrS+R27WxjYShvGNZDWTKANt2ZR1o4+aVtmEWX0RDI+t8S9KRHru8zABHc9Rqwg422j3f3NuNmBeb5NmNCLsdHN6T2fPNwsq+LjyPYf4m6lj5v1EVm3/dcFfcKffyDvNtwuI6HT+Ye9WBt2nd5eBJNGZlTipr7d+bYpf8adordG91K+/z+4wVOtZfehwC1OVtg1fnYSx4YGuxHI6yAABHv8XHvSCCkpM5Em4ykXcUVhYpZzsfCDVmc2CNdILFFbppZCk+cFI5t7D5KCc/rm0r/azrvjgHeGqS19mD3zq7lnoXlz/3KXTEvjyUoyUP2IMrPjwvifxgIdErgbQhXHAWweHiLcMUW72HwVAz+iHlg5RSHpmJN3jECIQMhDMuGR6BJHUBhf/6Ejb73O8KkucIaiTgc23OGhdaN9ejQftl9Lwi0zSM8TkAIK3FRjYNxhPNzcltHltlfQvkOTJzqMgx43+Xld0CeiS3nDbyHR5YdYIB6pEcWoA3EIDITHlwH5KVQjsplK5UhSdfRcuT8Gsqf1rxiMJogi4rhHnuVymUoTivk+TVflND3KrE6rYGx2BrJjk+Gu9Vy7IsOuQ9AxeYqkwZyVRnXZOIUBcaRs52fTCcH/bnW8rMSM2xysPguRMxxVupocVaO2QI7ULd+XU5U3kjbcEqhKg3ZZY/DHI+A292nIv2WzJzf+L3BHqzeZkykdYiFr5UntNn3ivV6MN0aTx13oa8bXeLTf0R/sz5KuyLiFd4AbQrMtkdz1qVP3bEYheM/UoIQrwZrqcERvIDEwroJrRIhjcFu16S+LjhZtpV9hJE85sjHE3JSlutpm6QSY4lKZtNlgTsjhLhyFY0bGXToXwaOPAzNuetsVZwVuiCR90L/G0EsMZhzcBcaGvJ3zkfbpuQuK3rGkj6fd9GORyz+2L3TxPk9s6EIgZyJMF9e75Lw4qOK5DIebdRPwuKuCp0AIHUS+JvpWIYGgAVn6rz1u7lM//MxIiwzsRvvmafEohUn4LE8DQZuDBOlnqUuJv7GOMW1+4+g1D+aZbMy1gMeVXSImBAPQuAbwc8tJ2WRngiAb6WifVTYo8qk8xte+9CSaeyTaucSXZnHNlB/tyqUZTrR+4S+R98Gm9E0EyA6nMr6EhCMqbhjd0mBLtE61DDYk46PbYZ2dUyvuQnHacIvRy3GXmfj7Q17xa9GwqFsU0TgSTdEVkEl3WJ8ata423CB6jT6/GTUHFXbg1n0r/xR6k44kmmDXOdzG0xh1IJvtS9wjZ5imGz6LEiKJ7zQEtVkNxt0xvpPxu/1xS/0sszjJ+KoqdAWT0VMb8eznoyz7JkMJwSuoKjf0POO0sR8BzwI05yDyog16i7GtbTJKiqyKlXfpUgEa/c77lsYek+c34rMQY34ZbsF0rbc43CEHRO+1tY1AwozIuCmyO+axQzJDiDHqasNS0LLLtWz35xSoHJc/H26n8LLXRyB5F5mS0sCKzE9jeiUGZE9UNmZ2PpwuG4+bxdMW3DK8U/2gGlGZeRVOxWOn+0R3Y4ExwL3NvBU3BErSCbcXLAp63PCJCp9idy4jyo7W4YXxwQVquH788JaDFNtkUKcudmTLvS2cqwMg8/KMlEby//wwxMCalwTSdnZiaNlbqbHVBXEyfmMKSDFLJdV+hGrA0ixZwGVjZIeLDKjEHVFMmVLfitspS7R+KeORyGYZTxE9CLdhJcUQjK3GmS+TsbXKQKZ+W3CTrNtx82PZcEHBcBczOG5PkJiNQdon3BGQVDupRenAymhnPLfCMrIxMG6TQXMnKyUkWXf0DqIdd3Tfvg4iW/xn3BoAPG6TF68ZCoXjYcz8t+FNpFqAduxRGQiuPIRlvrosAdB1MCgy2fFwZ720p071G8owUSx9loDHbz4dMcOhQ2LAfMLWbOgBZbZ65EKZwf1z+uSABftJ3tv6teipb0njGQvy9EEdFfScw+QwihC8YiYKfaTVYFMML1IzVQtux8j0zfj5OR1JcSOcEXvclTO+Ju7SGVk77jkMirhNOjN6iojmKDxud3w83I6mdCwWhVW9xC16Amx378IJq0MF4W6Rd9vHrT9h3BQwGsEsap8628hBshEQvd4ovTHCHE/LhABf19qu8CLLVA837bsBO1TowriXD9qUiY6nMxHsKqI+02HnzC+EvMlpRDnXbM7JshFJL41WYlQVrGEeShAtXlFFIfg4p7DERGKoG7KMhzuIt2fmFoYjDiB63OyUPJ1tdhKpis4KxPcXSi+/3YsxCqWMdIzaU4rc8C3t0SnRh8e4uh5ChQ7rp6SNmBeqlqlwl1kILznAsOHkP8XZO2PLcuEsl4eqel2bLnIQy7qifZa44dqwa5jtfD6471Bu8VDK190XfVuaQbENkS7SGhlbvmC4ZeNezXSL4bpk0bHALZ/iXacWmS2VEaWtfaT03MreXuZrrSLbiLplJHaLlzIj+cUnemvhuTV6iMLkPvWeaNcDpKQBqWDqx8nR3ZP7c7gFE6/2FFqEubkJNVB7k5nDrQKktkTYNHXHzo4aN16RQ+Thhl0azUFIf/q3OWSTqzjlLNP8uLwFoBrQI6L05CAAGvLRWge9iw2bMTAvGGchD+YDDfFiI9IDkpLb9WUbLPMCd6Q6jd4v/IDHLUPYulZn6Aqq6sDMKdg1bcGv5A391uALc5aqDzAeopycyE5A9DnagjAvb8YMs62YZnH81KkjlpkrUb1ojH6rN2JvLqCysZjdc5Rko8t/16XwuZgX7H5uSw0S7lpbqEWM54dtG7jZMFtwC180kprieroqoaCFVpigWRFcNuKdXWvRj6kv5diYwmtTzMIBo8BeMkmr5TXRC1JkQJ4odoueGrhLupm20kEUWYc7Xm7LGAo+geRXfsSAStyOOmpXZJRxS4aT+RpkX1Mnb2qH6AiA8VD1ihcGCg65gTOJfD6W+sEZRwuEBm4+6Z1KWzEfiOgCiLYJB0UYApqe7EOT8TRm8plXwbQ8JGldXispkti50+dMR051bXGMIwJmPCT4rKiyfbvbvzO37XGXdBXpKJ/nsWKp3A4j0efap+t0KOOjj7eRoEhddCwjGOG2TKesiJPiG5FN3E4Zc+TX7Kyg1d1P9LNOFbhFrG7KtPjocCfCGabyjBWecbvmQkvbWd+iPDhH7Za4qTDZHPowbtHRki9AG26EQEEx2Ht6AhBA2ZJzxMXb2tqcrNNnkQPsmmxo4+P2fSKk3b4jAropEgSNCJGWdGsXkcdrJSOkTTEsET/PqxfCYsHnXqOCsLecJwW1abrmhsLiaHjeOPXudioP/g5OFRV3Oe5EGa1ZKSzKCe5ypsdwl0KB/c2RxPVDuBELOoxvQelm3Pm9UbnewKKKMdqq2aqTA15dKBRsrOsyHXFg3khsPY6nzX+azqMxJOH7xRe4NLtouzCKoJlUlcbixE2HW9PqFprbcJe6movEzXVIxCceXo2Hu6xZRLtftu5T8nK/TZp5Y2SRdzTagsxewXCjbKN0OKVtyzM7iN16bBRV1YPmpzDmRhrrhRzF+6MwMq3SCgVcPE1KDUnTouzTyQYU/bLizOg01ShvTGrSlBwOtV1E51iP2vlQ4iq8dYnb6WzOYFKnxS2FM1DygkUWqm/Yp7K2AitRUuKQHWkELVHPTIi6LgLQIWHikuEWZW3QRRgbNaOCH7ElAxFZy32BsjfXX1MnrIsSN3zdBzUANvxkIIk13D7jRjtu7Z+wFUHMYxcH6Xe20jVIIusAj7uo3fi+pV9f+0l6Tc87uUWOluHYzFBUvokmJDvJbTZkTBhb+ubvRHpAFaoQ/KPIuajlvGZuKnjB2nseohLnxmZ5jBt4rOUiNDPLBOyjWIDVPfL5qmNM1MuKtqmtUHXsb5dCZwWIz4/brjXlcMt2GXcV5NVN4MeZ/VoAwZvbLesuyLxwfAOqqkuRJPh7Qyiuz9G2dZhDUUVlVyzySi0UuEG4x6sXyH0kDyZ5HOfsZskcFqRsiXAHxOKdJ5XjV5I34W5kiKyvLbgD8yZf7ZyDry8035UTXHto1anCDlpsJWWJ/vrQhjt/q567gij3SzU2hyG3rwEu00zyDgGhG0IoOQUnPE0Nm8auL9nNBOpQhSripWLoOFR8nizAEkaLYBu8lelZ+2aPKT4/HQrEMEk55XrGQ9NDDdzMw3TOpXYN3Nmzs/cXpit8wS0Rt3KQU7M+8vl6hWG0jZWFh7wLU6Iv6hRkGVHZQZOROtroeQ/JEkRujJvGtt7hS0/RiI/cXjb77DQ1AkL6St/q1tToRccA2eTWZy+caZY0ed6Whi3666YcFTf8dYV+mu7zCevPZWHKKy8OhPyGO86qCmcXRd6ICIo1OQAd4iiPacGW8pcDsXfUbvRANZZMY6x0R6TSGQRpJK83iGPOu7rIrkKKuoGHCj8CnKpawbHlo46itmspCtibq+SwnMuOUByFSKCUaCOtFNwUxULhMHK/unqQPTHhjjWl/6IMJe7yo44iX1cLbnvXpGQxyY9EUwQyQjFqh9alvUV0cQ7CoqMs2lK+R+uj+exGpqeMzLGoLRXRTcfQqhfSj7xT1dqQlZ9+OTJ/xSZuh1kMkpycMJ7knQJVxk1T4EGcVsHDyJGZDY30tznLCKNFcNei12N6n8q8gduci2ii78J7Hr/cvJypkQxGglXt9NNswPExdEOogosQMc0npwU5hbdRbkmhRICLN5NimUTtDKKcWqSxMIkAPsoXHjbWaWfuIn3y4zpqh49pWslRpPICVoPmaV92DCliR4xlHtlKvObYUomGU1KK0s1iFeOuqIkalW4gFAGZI2exFLhTazTsckPDjldkkmVznw6Yo1JZ58wlyPZx48zISN+WRuRTZaQzDJqpZrpCZbMCbrirtQnGTVkEZT26jL3kuQ4xQpZnE7fqTiFHL28LWIlLUkuD0aW8Zb4bfB94qSbhcMPfm4NdIi825Cz9l7jVAQtGDn4alEvc6ZouEJySJCOoqDtDpumXPsgkXjlnEHk/SRvBZG/YNtVWKpbrkc5lZuvDMUUbjQ1olKE0S+CMpRhr0zjAvYFJhBQq6ztUukTcPSMhytIYwpRTqxk3jzti9KtUHW4U+Kj9si9qOzojjOCUP/L9PKyKtJUe4fb7XXD2GbVthytnJ22kNXkhuCLSAjJyLG1jf0dDaUC8WC4ZkMYmwGROwyDjT5WempWrQ4A+LKczc4wbHrc6Eh6yRKJHftN9XBdxw5LgWsnEj4M7tjoKW5EJr+tg28wPQlK/nufSpzjIiC537jbl0BtsRiG61YvBgGRFaN9FmNMZYrbzetETrcxmjlGGgvKSlnu1Pa9U+lCVyrToR4RIq1GjDFNEaIKTnYyjlbCyhpBx+inW4hr34ap6oXSNWRTrw+EWltuPFtzCR6FDcAsP2XAzbp2e5jb8NXo2ALbhTWFQfDnJ0W/HyA6wLjAm/oTKPzdigbNwzi6sOwLRWH3s+Cu4K2qi4ItzoLBAw1PURJNvpgU3aGp+HNxJL2q6n/WPaRS7DUhPE5PMGLe7R2mNVnVpjQbE2Gw8bizTNi5Wpke6TuoUcg0gwxRbYVnlsZIcq1RQNoaiaBsoAqki0XCnEZmCtRNCO14PXulKuPkUzR61CqQddxDnyhlRiVucEaSOYM3bebs3tc1RsXAewi/lG+MjuohP4+JGG24+R7j1OmQblb68DNtxF/KW1ZHqyAtn6HhiBMvaC5utaLBGaS8fqAxq0PzPY2rFTY5AhgiBcVeCmeSbsYoeeNxCfwtu4Ul0BOn1tpaIsYrdFs5EZdGGO3XQhQqmjM5Q4VmjMjUGI1KHIdG+HVODozbkim+iOT/27KIGgEDGFKHeOpGZGanCL+kTodv6e0tAaqNfuVgau/zO56LwoTByvQbFfTHRKMpOxpEUJ2qKrGmgZgv8zAA0khiZOUFlRxijPXSWnZE+KETtmJ21G00gWj0eYVXI/CXDdTUAlof9TrUhKuCJvsVIMnw+3GJIApCivovwuY1gRVF1drGGzdwxrXBtql5LpsIOpjElmXHbBQVueaw/6n1Op9U3CV3Ph7vM8CrrUmSHLG8ORrHWxWimN9wUD5NtBMG4daat6sQu7LFBmOFFi4itjoB6LFJoK6Dw/gzeKAMiLfUl1EpGUIHLk3KIdVp16Lx4Wy2EF5jQLARhKGmzKUeBThv9SPon1LKiEPNbcTtnZMfE3dk1WRchuLNzQRvu6HGrXKKJMtoOXPYwkBRlBXcxrRay82YHJhEyt5muGaNrQO0CgCg+484t6DHDzZvVmIhoP4aKaGzBna4UXRU55UlFwiLTjOnC5FAcfZzeN1Q849HZLhlqc5HbG28rbh6iKwtK3JwhgnCTDQIIeWPtRGuFqNlNi7wlo6vKgn5pz7xqFXouRnn3TR26ST1tbl4r/BlFALLQAuTxZ+tPpmCs0yTCNJui+1bk76TAMvxocRTOqZinT99U3XdZEAPmqA7NXKAYeEG6MYj3GBDF0jSYFF+FSgpefoK0b/4TwmNOMZvYKUZpdCpx19CdpfXqaF9BHCRt4iIzKSEQbpFDdh6KSZTWp8O2hiOicpmJyJroz3zTAqMYbSMKC9agytk6XNLhgV/To46s4bBD1ssSt+iJZJdBjEAdF0huiEEdf/JTHNDkaWJtKd9nx23GxDtI9wkAasZdXF/iRhvu6HAjdGCzVOQUc/AX3jZmvvR9xAKRZxPTz266oVN4PVHUvBIu0gt34Bfj+MiQGBT0uQaYlwpspEwVR7FgXpSzGkd0y3oFx9yo/WVW5itMEa2WyrM6IOYZbufRYUw24wRkEZpFP4lSLbM1RQEMopC5HWJagVGm8oqILcRoNAHJJy8nU/kIPWJwhLuyY8HxOHjcTJ8MebTwGzS6+xpA06FB+O9wG0+avy2TkeDDmYBQnqIpnANwhluwVeslMfPYTkAyZcMstFMw0X+1yTvC88XJPGc3gpsdKV+nv72DiIw7mIPkOTCt0bB8IA4y/3JD2Vp/ymJK70ySbLuhqmLg18U5wUhDKaqxClvkoTltTbmsjYCQg30AG56JwHt9IyOqEZoBUEU5e9v0Z60MiLR7VHKi8tZ0A68RMAT4h9xIISMA3azFHJs5PNED6a+2FDpnaE3c+qQC3MavjbUZhFvwRTovwzRWoromhxzzmhSbUw8SYRV3KW8aTlSBjEQcvcibbpd0XlN46k+u56wyiK6IitTGdRprt+Imnui4Omc2DreuZiUfJtOg6hQYetKzKPqTW9WhKOm4OGNGmGSZj2Y+qdxzOxYDxaBrIyNaph01cNpQQh8MQ40YbQgrQ5Yq65ziVnln3FXpJIkB2VlZWGnHLbrQVY+WibSomxvMaVAQD13xw0v5PHlujWiV92iRBGykcGfytF2+Qzyc9mZOgB2Gc/wRmj4lOnj5LDkF6ZPG3erY5Zy+2wNIG5vwgiFAshLx3BFQ58Xd2DBEkZm4lGc8XqxUeckdsG6S0iIJO+OWqJMedJIIA3NM3AbhFt238bcYW21Zp+NhVPn4KGX8jBp9c9tRphBBusK4xRhL3OKIoLoFxLzcv4kbJG/uP9EVtF/boCdfSwW+pDPmdLigKHYwPm7StBBs/6FobfImNaIkile/TeZuUZXINAeDdMZmkQAzfFVAeNwq95xlag0k42YeKD9DlddZ0COxIqoQbas7/5ap2jNLDVzGTrY+we6haZx8qAatgsuOgrOMVNxMmYJLaRUoGS9vVYYqK6c4ACtyNir+uRBoTizNNae3to+HWxhKS5OFoWXYihLhhfS0AjRkGtMlVFfJfEzeno5Lei8pc1Zq7/Tyrub6d4SNuzO+HHJiHDV+5CgV5FrAtgiIQFqxKmTwDlhZXiHTTNgDIuyR8By8nbyjBRIOhRBDyrgoPdAtEHSoJ/EwgNef2ObD3J/JUD2j0KzBpqYnkZECV3ZeWnsDTC46HLTvACC9rjNatqe6AaTsnB0KOXDlIeMWJ9V0wn4GMRpuF9BbcNPK0IRjTNemBAnYkfRZdWYsb6uX9zYQj8cZQHIKHSI6eOPV7fRgyioMElnofpzCUhSC5LGvdyqhCtC0mxVFxnsulAszrGZiU36sJBaV1O0DCJpF/bO4JSrJeR+sOZ2Xh7rcTEndotDGdR+ZeHyvuCly8gItyRJg33pcI6U4R8Id8x3ytKMoqYVKcmB+diexMfO24tklL28bMnFbkdoMxEDLJmObvFFE5EDZhb8wO5ukGyYvmoYNAUG3amDcZuie5uDIFLp1eXq+hgjIGyxXBWVynemP4aYl5/mYTMWya07/l4ywUzQtuIv8NpL+6qyT6J3gNmcWQt78xgKUMSMiopKNVKKIxQxJDDMGMxYBntbVk3Hw+FiUVbydVpZDfrSbHYtFukjC5fgtQxwG5VJmLaTKsUKJ6PVG0naouo6GdJ14/cyS4JmfyNYwBZ5etMxDnBk5HbNgPdeO2+ohiiNacdRwqzCJ33L8/zX2plF2Vde56DfXPtVXqTr1qAMJ0QmDRSsQAmPRhc42mDgGOzaxE6dz7nh2Rt5LM9LcN+5I8l6Sm8a+17Ex8XUbA8bYxg0GYywBkugkIRAI1KOuVFWSqm/O2ev9WLNbp2TfVx64Sufsvfaa/Tfnmmtt5/QkamZ0B2WuydstCyrdOQ+zFFMd9mnoVgcuaZEvcDr6SlZuno+Xr0xEDxP2NAvd2bX2Y70ulH8fjB+op1tolMgrz4ymn6elmz+zJVxkztx0QVhepnob061Lo6ejm6Ib09uM14FfTrcu75M5daG8XraetxXEGsWYzodIz+FbIpIzkEv95MQZkFc1B8d8iEXpmCMFk5pT4jJ/LqAnHYnvtpOK5RHR1URSumKM42c6wSvBugYNJ0j29BJdPN1ZIKunW6wnKi0z6VZVgtQ+DG57RZAiluNfPd2CRJxBJyX36ORX0K0OSprC6l7sFJE5GJs57P6MbuN3mm403ZBHgXK6lRYZ2wrBohtMmDppnYuvMWggMv5BZSh0nIbPmg67+cfopmVIBhA+EXwo8afmZSfouf4G6cTM+lYyo+e5kX0CDUeOp+qE8ofaUEK30+uscG388S0Oqu/Rj+VsWRG88QIAKuIdLUKT3uz5bJ8leK7eiQUT6xTIR8DEmsgGKizx3r1+6YfzvkSm/n9GfuQ3Y2lR1l8hSi5/e+Vwv///0h0BPYcUyOlWgfmbSK/Ldk1qdPLR3W4j7omg0/BEz2sUR1faOr/NM6dB6RYFFaOUf3ubqmewUkKAyCPwGr4eXVenyOpQoMYuq1PJKZyGbqJUH6O6yJedDm/zPi0ycEfSZUgyOsKyvx2PiGaSzmdzJjXJ0bGtWJhRKm0yFVew1DqZRne5yRXGZToOfVnsZT2T3okMTdgM0t9s5JH7caR2pQiOUM+6jBLWc2eIamcRlF4ypN1j6shyLTLhE+RofG1n5esljdClRsojjr6BKROieLFoCiT5s9QJxJCVibGuYSRYXq/j5cJMhEd7bma4vItUHZlTAPUoslRlqwBKN5lhM7fd46NGRTdhjiFl9pnc5KNlUjS3khGN76EwxxI93QJfVXFi3XNERWo2L/oldMOxK6R70iwNzUSRiYdh0dFNv4Ju970ZrETBpGtJYU0vA52ObhY9nCPR4rTUsJzOzdCP3MGJ3zN+2JxtJcf9W0gXugvXt6R2VOoTrG5l9wFSO6A09yB0E+u8HC0gxNa1EajxSlCRIrWTrX9vi+oXQRc4NJay045+zpDTvV0jEQj5i1D4QRLRhAAVvo9mZPDJ5KDfS7tplmfq7ckIbAWCMYUULCFMARB9CmHCtL0gHJm0cFPHSD8WrCOS6lACOceSHIMcc5/hASPVr+6oMABbRakL4/yMmQcCOSPI2teBsqw5/sGUj5+Nbt+oAAAgAElEQVSjTUZyjxaX2Z0q/ytuBNfzgdPRnUN3qjuAOau+u6htS5OOqTPo9jzx8snpzt5C5ukWZQ4usMA7/3q6Zcw6hBCh91jqwEVDtfuQ3a8rPjohno+gPsp1RGsd0VCi1id0EPmT3ZcgMyGFEt2KXdyp4GpPRLq1XpFRvW17eVNxWv6oSyFCCcQKedXzHY1A/u4JzXXJyHcOwhphJGo7T0/Ws6B9BAyrfCuxAUJe9w0p+psxSG4fEagCTaGcsnoztkN34I5dN+eRCdTD1Ky119PtkULMlcvsgOcnDoqVhMQ4JBI6R+zoViUlK/AZbanoLHzI6I7mnDI4W9Z0Vonc09CttuOcsqNNl/sETZBz+uRu97zL6HaniMmV3igzJEOgbPVKBiv0k1zeTLfqLetIWXNjREe3G9s5Fw7x5mRm0B1noCgC3P45Y4QghLQE7Uh3MlC61S5Yzz1CZD01PXf2GAXlsnwd+jIELQHVHF+eqpIby6Tg6dYGNfB7Q9QrwU/UeUBYrmnNIKV5VWWWOZK81y1CIr5AHql76D3qYRNBlC23lhxorBnHjy/XkVcWnmO2qw+OQcowOMNleFlPN8yRJRp8LwDU8wuVsFko3eSWELWirrS4ZUZyXIuOx5LuaAU9OhuzyJX6SqKdrqVK4aKbcc6Zk9CVO21Nu+CMXgyDrUVkICChvpPVJON4mqV98q1oiyAtRmR6UphLPU77E0EoEH1RXZ6f0W28y4+T842ExqFMlyRyyxBCN1OZPvOrOVFMz5wtvEwNVSg/tD9Dlj1zPZcJRnevFIBz9DOT7uQErLHMZOw1VuYjwTYRXVHj9LBNHIP2PDg4GiU9AHtfhwoi1DOa24ATgBlIyq2dMWukgQmazJmYIdcrfOa6eWiJJP7N3vLbQz5pF/dRpqyjm7v9pCfC1ykc3TmMs25AT7e+cDmLHk5Jyd2rY5V5RINbFaijOT0mmN83i/YXuigTMznpPGGoItFtgcS+Q3JuPJfk51LBGa4t2VCCl7HRrbtYvSMndqC6i9YUub4cqbxwqOiX0W2NXVCDV81QaM+OTehifZOCq4hQaIn6XR3d5NMLiQFeH9w3mvZ4I4Zem9ViYIFCkbqO4x1FHd3Kc3K6Adhiguh86UCNNKglRlUkSuTeGM7rcSSURhthnnoym4D+rdGExxZo5I3cTUaEhQwlEfsTy9ENhnlPLcUmvi/Gun74mRE0kRn0395I/cEhfpWEyNMt88cMuq1i7c5xUJ46gdXRLb52Bt0kfDTHGEL9+1KEp67wC4loFinzSSeiJEgERTx+mToy3XaatI7lUKRE0DRPf8YnI4EZdNtz9YAXJESR8n1DHzZ/d49R4GhiA3f8sHzdzcXTLftNfLFQ6IYhAxNQnobPpNsM3ej2Zu5pIJN36buixdmb7gVntPb0cgbddnaudJnW67jQHevmKSxLz7SzbjWUIgKxQtIgJUbimQroxeKNIkkOY8K3vJ01XhgNUXr2vIAaUe79Hfwj/3lqlxaFqF9W1NzdzRbusNRIJQh1XZkOOeWvKpAKO1RBsloCmRCIGT+DbnEmPHfifTMyH5ujIJbCeEH2NEK0vFznKn+aqD3dVqQWpZBORX+R1ItKnWdqp+f5Kd0yC6hymZKizgjTc4M2EsmmJt/z4QKQ70fgOWkkB+rotoY5Sz/8TBzdYgyuWGvBmx23IApAN96px3WGOBNVmU34YCAORRC5X1LP6PZosY5uOZgoO+QX0TalwfeB2BXZUQXEx0GUyBE105DYQypv/+9c66TeY8jVsuACFSBSqupaMZDqVx+cL7d6gDzIFfi0eQfQdWH1ND6akmNOrFMsee5pqrMuss+Emk44mgr5JdaM1ex/6hp9fPqk03UxLDpkIsoh9PHz1QEJqvHwA6LcMg9TxoyWOocJAtcg8iJx7i5sDtbG7Om2scSJkTyLuCHP7dj1m+R8LEp24ldPGLk5xxszeed0K85zX+e1FT9XypZK1dnU0x3r6HbPzXRJHK/8W5BBrKM7mF5k/T8Z3bku6LMkMGrKKqhAOpbBcxWHdXo9Dpme2+dZuUB8hfA4OMTvPstY7uiuR/v55jqrb4AIsVZKZ0g0yB0Tw3TrrI9WrNSp25MNRYwh86iiQDMjgV4bY2pnjtHpjiiDw+UuOIqjArzBOmaQf748x3UPOuVRZnksL3QL9K+jG0q3E3CWC0Qdh0BYe+0cfOa++epU5XyMlJ74ZUIo3cn3eH5yZPPFwKxrM68DKM3aSWnIMPvemArEmm4es2gsqQBY3s6ZKu/kYinQltmwyK4Vut19qmv4pXRnepjRjZwuOLp5rNPyxc+tLGeMKXSLnPW3jGETd3865EpubA6E9h4Ym6tvszZemt5JyqFa6OpMxkP5u9QxfG1Nx9W0kgcs0ya5QPW7pI1eQSuC6AhAJb0KkKOsUu9YSnVCiQ6aRf+F/W2FTPF+zMroliHJRVnxtpFXOwQGSoRyiEWE4pdq07Xp+QSyU7GcIiRY59BHSC9gDoGr545l2bO8MrLQYlln6I7ZnmldTcAXHurj26NTPLdExjzyeaQ+TyOHyUOjWXRpE2zsRLeLaD6yAnpylsYyw5mObsocqcLTTNaOJ6orycELNKfooxOQIVZyqx5UN2Z9xISspDGtQpfWc6A81DSQoDwmIMk7c7j5g31qqQYJH6B89JdvCP6Mk+CfQUCOGmU+0Gd4h68BjenOV/vsifqbADvOAPnKiyBQR19U+RjdIhtCRP6uH8c+R3GgsiRRFDNyqAOBY179kp8wRKOO/O3lrl4v1jHALc3w36KU2hXnHIconMyBlOnihdmBuWifN2mZ0GROpsT1dNNMuiG0ydgkF9t3AtmQUNPjTxzH6CQXr3juiCXa2grMn90AqR8YTQ6tESuiRzGs+LI86p1ARnewuomJ3tHt6LWYQBndQjkJrXKp3ufkrRAfaG8PmNtdQLb/d3c3oKezsOjH/LRGNTi6ha8+BQXItS6b8wvOySKj2ys4Cd2A8dghBHkfrBowTJ/UOJ1eC58sazLextIhm1+i/4oYlG9ODCJ7bwdCd7aMCSdf0rTJ/0ipQMbURQhHdwo6Ts8jHN3kZMPOUBqfhCmBAkIoQKFg5yWbzAJX4Y1hgT+XTUlEga8nZUgaK4BC4LGDeWIHgzLhcDOS3O8ZKLmcVNJNkAbbSAw42DxVes7BicIRhRl0hxl0mwDtO3MUyi9+fsusFjz85Ytw1fmtCKFgWhN9qy/rxafumpvxUvgv8DBdb3wQxUk9FJwOSYSMjm6+VuZKp6M7GP8DFSqjltYKPnbvEnz1X1fhew9chG/+ywX4w/sWoqutouMGCo7vhSqdKPvlV83Fb90xR6+9+ZaFeP+6LlY+czrewRIRikrAf/u/VqCj0dEdpBlP+i2CjiEKLnqjtEEcuNAtnwczgxBML5lHRSg05w+MTCkQzyE43pLZhKM7FBUdT+QnMq2n24JMoiO48QBznrKtQOkmR7fXPdTRLffI8/j7EJI9BbFRIrXNZLuU0W06zjzTZRuenD+dSoxU/8erJmXMT7DSOBRlLEMB4lmz6MrKm9Kp0jwfIrTZi6yliTVFn6QRyM+7fp4w7+oLbgIry7KmntfuN7pnjEeEUmjx80Lp6IaCgGvW9uCdA+O4ff1sU3gCsjM0kybomInuYOOTzUW0LRW4hJelXaeyEONydHMYjDGijHzYCUjpBgFtsxrx//7l2Wgvp/FHf/YG7vzEdvzB3+zGeKUR//inZ6K92cmD8/901JvN7XQ8f+aZY3hiyzBAjsNe8SWih4DlZ7aikEUdD5mVryZXWzq0VMm3dxvdMLqF3uhQMl9bxpL9rs09lmU2fhpLxsl/Uv3NPi9lb4bqT9LhjG7yeh1VTk7Y6bfSLUVS4U1uf4p6OYhExKSzqse5LYBki0WO0ISPNnair4IQxP6Qtfs6OJrGNULSs0pAvDVJc4owR2BOdE2JBvNUkBHWUq4RXviYDEdciDAwGbtMxfVE8DMkwmrBkKyxSpTUo5EUFng5TBqBhG7RU/+2bshu15xubXoBgYqA267rxj//0x589jNnYWFnwOGT5vTE/RMRGiqp4j85Hd38A0IR0FAAE1PpeZUGwuyuCiYmajg5nArDkvM2NxEmJlOe2tgATEyWTGNET3cTQowYPFVDNbpUwwQJxIhPfPQMvLb5OP7HI32JK0Q4MTiFB76yH4N3zEd3e8DIBHffFgGzOipoaw4YODGFyWlL00RPksxLDPRPKcoBo6KuzgqaGggDJ6YxVU10t7UUCADaWiuYRA2TU6q5aGws0NvVhLGxKk6NVC0/d+lER3uBjpaAgRPTaT6K1gJKPf/ByQDRGSHUiOvTPk3bQPAoXLRSv5OzMnlMa/cPkPfBaO1D9nOoPfAep+j2/Widzhyi6BmpXUqnK48bc7qtvihO19Md1e7ETlThnS0pCioKVFCWhIpjkP5Qdi/EKACkjk8r5uhviMcO5pkZIXivqZA6exGQGHbUVm/NyhhyWyR0HtdBdF2yAqkdpOclqC41A8hzdBxzRp5owSJw11nH6Wno5s1ry89tR+34GPb2TeKnm4Zw8zU9+PIPBkwRVAYBZ6/qwqdumoU/+rv9uqQVEXHTLfOxrKnEF743gA9/YD4uWtGMvoFpzJ7ThMmTE/j7L76D4QmgaCrwpb9dgT/9h3343Y8txqyyij/4b3uxbHkb/svHF6GZIspAiJNV/MsDB7DzwKSSJMGto7cZ6y5oxse/uMcO9WG+RpR49HtHNZAsO6sdH797HqhaYnQyYvmSJjzy6FE8sWUEsazCmJeu/8Ddi9A+Mo4vPz6Izt4mfPaTi1CbqGJsKmLh3EZs3DCAR58dxp/90TJ0tBb4k0+fif17R/FPXzsKALjl5rm4fW0XjhybxKyuBowMTuJfv3IYgyM1UIxo7WjA7398MVYta8KJ4Rp6ZhV46DuH8f0NJ1lXrV06cwQg1VUtE3OkJ5J9HSb3iJiOHmSUmC7l5X/V8+gCLj+v7plqmA6JiWOSQ5fEqRAX4c0GxL9bUVVVyjnOGO3ckwjn7BQlAXayFn+a0R1sTHVGQIWCz+kd5OXQap5JmrY81J35o763LJ3BipfmscTIowlTi5mIuvyjnk0YEaU9XLyuNX7J08GoxJpahNHinaVjj1QAEI+tj6IUGXRMYZrNt/5HI0lZ4vb1c/D4k0dAAJ7eMIj//tnF+MaPBjBZY6VQtkS88eoQGj+yAGfNKbC7rwoiQigK3LimE//9H3cj1kq8vuMkvvHtUfBBSvitjy/Fb97Wi397qA8xEkIl4BP3zMfXv34QO/dNoHtuE/7v/7IUn/vCfjy/YxRAxMWre/AXn1mOP/nrt3DoRE15HmPEypUdeGfPKIYmkemC0h0jUpNJibJaxee/uA/HTqRzPHvmtOBf/3I5drz5Jg6dYGMwVTZaAdz9vnnYtuk4Hn5mCIgRRYVwzrJmVMen8Od/txf/61/OwV/93W6cnEzMXn/jPFy9ogGf+etdmJhOY1x51Wz8xe8vwh///T6UgfAnf3Qmjr5xEp/8/F5M14Ce2Y34mz9ejtpUiR9uGWbV8ysPXt5WE9K5+vTH9yuIHkv2kCEVIFtp84FXPLIEp+g7oR0yAWxPiA7h7ADmRNI0uSBJprtQNGHHKOTH7KVnB3L0e2eidmZn8jqvhuAbi6ReIMUOLTAlSvheK4xAGOjyQyme6aYWJQKQfbaWVviGLhtHm188PJAGJu+AdAwpWJEHMLmQ4RpoKBWpEm1Mt37uaQPSeRcyNTe3+vlx6tPW1YCLFxfYuGMMoICh/nG82R+x5oJWN2eeGSVH9+ONJ3Hzuh7l3VnndGB6YBz7B6soyxpeft0cBWLE05tO4sJz2zldKdDYUuCR7xzGa3vHUYsRd9wyD8//oh/P7xhR6l95eRA/enEUd93Yq5RJLt3aXGB0zL1bgxLdV6/txd989kz8zWeX46O3zkYk4MCBcRw7WVMSTgxM4vV3pnHO0ibjmwSY7AzPiPa2Ao2NsgsSqNUiXt89PkNmAEAVwodu6cEXvn4EE1WdMTY934++sgGXn9uKlRd0YUlLiS892oepWpLk4MA0/vE/DuG+u+anhVrRPwvBZkjgYi+ZvskpbmJ8M1fAolqzHccvKa7R7WtzXj+Q6REy20mzK+s+88gj6H9abxPdrmvR1mBINoYiDoD1n9w4buuGZAbmGQEAFSJK21+CdAXWw3MjLLVuF2rssjqiKENf5Erm0SRF8MzUZzCTS0k45FeeyiTvKYTwfcpKEUKqogusUk+vc7PTwCnz0DNbeSMzP6lEcC3rjLFCxSCug5pEAe+9bg6mJ0t85IMLVcFbK8Bt62fjmVfH9Fp1kCA89cwAPvenS/HAd49jqgy45bpe/OipY6zMBW64fg6uelcbJiZL1GoRDS0VNMrZsiDEqRoO9JU8r4hzV7The18/zjwMejjr1tdG8bs3zzKFYMh59PgUFs7vSDzTFa+Al146gTdfH8b8pW348Np2FEUDunsbcN/75qKzJWByKqKMwFnzG/BSY2ERV3iZpV0B//nIUXzqwwvwr2tn4823x7D5lZN4+fVRVGu2giO6MaurGXO7Kvjt+5ck9VDuExbNb8DBxS2Y09aKHa+PwpXegBixd9coKnNa0dsSMDBpkVHrY0y3psOImlIQCvh6EETeZTXTERAhoIAYp2IooVsRs1wPlGWElIn5S2jBWmOPnIlraNgnDzKvIHU6oY1X0QQZCS+ZAEiabrae6A6hgQGCKyHws0Io0r4VlkkFMZLfIAbyezDM4CITp+cEkHsJjhRStIAjjiddn28Ac/AMyMZTGMjJDkVoMcvn+1rJlqKiji/VaBFCdAKJiLGW2ocZ4kWBlYxYhG7NYd3adlRHKnSnSrMUkkABVAm49bpufP87h3B0iM/rQMTO3eP4g4+fgaW9BfYP1BKJpTnm0ROTeOVAFWtWtWHznmmsOqPAA6+PA4i49j3zcOWKCv723w5gcjrBw7PO78Sf3ZOQiLVlmROenCzR0lxotImICCC0thSYnEz8jg7y7tk1hOmOM/CuZU3Yvn9KlXdygjAxPomWnsY0dgD+6jNn4stf3I1te6ZQliWKSgV/8pkVEIxmqyMe1iZ5Hz08hr/6f95CW1sF557djuuvn4d7by3x2b/fr6mk1EmmqxHTkzX8jwcPYXhSTn2SyEmYno64dn0jWrpNbyRyVpob0IgSUzUx5aiyFT1O6W7VYL6sAESpndl8wB2YsjszxpKNTFYahGQXZBUtM3ItrT/IBzstQvL1uncp+7HeEYIgQnaujC5k6dRqLeDAx0V7tS2f5hNkNU/RUkZ3cjAix2DrqZar6uQVVpnnTzCoMFSB5HkV9sinkg+JFyttE1gIFU0DfC+DnBeg69i+n8FBt8BFTIWJ6mLlb3EZMKfhGKrM4MjtnYoperomUKERXv6T8UOQ8w2Swq26qBPh5Dh+sPEUXtg2jC1bT2HLK6ew5eUhPPXiCG65thd2zH5CXxQqIAr40dMncPN1vVizpgcvbjmJyTKhgvNXtuKlrSOYrMp5CoTmxkLZbPrEShsjtmwbxg3X9pgzJQIC4aZ13diyLaUmfu0+Vks88O0+fPqTizG3s4D0T4AILW2N+MSvLwCB0NjRgIXNJbbvmYZEuRiB5ibmpfI15ruFWXaBdWRsLOKVV0fxD/+2H61ndGBBV4OD5UkfJkaq2Hm0htUrmzE2HjE6VmJ0rMTENGHFkiZMVyO27RjBhRd3oqfNR1Ng3dpO7N85hJGqbaVT5CA1oywVEJFIO7/oeMWCouooKY1WTGc7iZLicL9SUWG7kT6GQuG//zdR4Z5bUTvSPhTRSfUY1nTn949Eh2bEkVgPlIzjejbETkIBeTex0g2zE7b1GGKMUTyeQTHS3775RH0IoB7RPk+EBXe9KLEQLrkiYg0oqyCk3YokcCemCjf0uhKINYtY/F22rqz5p58TQarKsaylcUrrpJNKsMw18HtT2LlqBPBYxugWpyNOzJaPb3tvL3789IBFV6U74idPD2DdNd1oKWoYHY8477xZWL+2B2fOTztP3955Cs3zWvGh93biJxtOJh7FEi+/OoLbburFgu4CoYi46F2zcOuadjR3NmBWi8jJKQOAnz7Rh9DTgs/85jwsW9CApYua8enfWYK5YRrf33DKKVBQSb+wqR8PbRjBP/312bj/rnm4fk0Xfv3OefinvzgLu94YQQQwNTSFfWMF7r6+Gw2VgO6eJnz4gwswqyFi0fxGAMDoWA0XrurEe6/uwZK5FTMkiviLz56Fm67qTsukIeLyyztRGZ3AsaEqYglMloS7fq0Hd948G4u7CV/4yiF88NcX4rpL2tFQEHpnN+GPPrUYa85vBQD0vTOKRzYO479+ZikuPqcV8+Y04NYbe/Fbt/Xic18/YqsWzpHpEq/IkszBmdHbVnfBuZoCU9JZ1RdE0wkzWx1HdDKESkINUbo8/T6W0v1XU521LemmTwlF2FwF2UfRcXbUUFsldYJEhkQlABpqFzpEb/WREqypWLZi1Z8XlcYGBjgQLpg3Y3gDF6UgEN9GVY+rkF7yQsoQgnjpzBp5rFS4EeM0iCWpQv3hPM660xy0zZnHcKhEaVEBl/q53zFJymWCLiE5ftS33cr4leYGnL+0EY890Y/JmkXuNAdgeGgajR1NOHl8Arv2jqNWCVg6vwkH3hnHwHCKSIPDJYaPT+C518bU4Rw+NIGJEHDv++fjPVd2YmpkCl999BhCcwMO7hvH6FREd0cFr7w2jOmS1akEfrHpJBYsbsedN83GlRd1YPeuYfzb145gfNrVX5wMiQi7d49i49ZRnLGwGWcuasLocBUPfusIdh2aRgNKvLFvAi9sHcK6dbPxwVtm49ylLdj47Als2DaKzraAN/ZN4NixCRStjVg8rxH7D05gbDri5IkqDh6bwqu7xvHui2fhrlvm4OZruzGrkfDPDx7E0HhEWZZ4Y884zj6rBdNjVbyxZwLH+sbx3LZRXLe2Bx+8dQ4uOa8NL2wawMM/O6n59c6dQxiYAG5b34v1V3Uj1Er885cOYd+xKdU30TEFoa5xUKO4RGIQ/BvTdQVCHUqh/NJlfEUKtsEyiq24KG4oJz/AKLKhZvpJqT/D9N3NVfWQVM9BkZde+egDF1DVdvwigj6L9LFZYb/OvmOsTdP6Wz86GirNrTYoHJOjOTXnaVCWygwCOTZAcz71u8oUhq3+bdN6jUcfsoQpBR0ZM5zmGX45yWFymZcwSJtp5Dq515bGRFFMeDMuV1QjEer0dPNg6oCI18ut5pGcLf8b4rBcniveyfd1uGeocp2Wx4aqTCnq6a5XwlwO5sRFB6T4Vfgv7HuffkafghauFiEH9ogC1zkspU3+dmv9HBTqT54qYw2ausIFE3hjkKtzeYvj0KV0udLplemlFRtFthr0lP/8HRGPyXRz9M738nhavJ7DzduavurtIzLdJjfXfuD1nIht1XRF5wlk/DQeljpXORYBAMrqxHhFxs6MTmYOIH91HzNS4AwhFflE+Z2ntoNumSEERH3TuGeH8FiICVqo0m3z/lpzYzquODmvKHbaE5KwCNBqsPoHsiIl053tGgTsLWkUEUvJ++rpJhh7DJ0p3bEEBZujLkkpKnJOUbpJSeKC7+sQI5XmM1UBVlK+Qn2WLVNbtV5YIo4qPczm5BRKjLS0ArYU05Ru0REpWBNA2hzn6JE3vwkfBEZLjUMezDKfsfTI9Kv+EIHKYPToPOro1tU4YWqam5lJWafjnltmC4luOLrJ6TipXOVzXVmToCAvcFZ0AH2W2bJbcnUSj+CVrijHCATIsf6+ZpeCCBc/ZU4iy9PZkso7d6zSPW1t30AZS6r4040SfOGVEWMXBM4nD2neMj1IfssyqkcN+VmRUQtArssyimc26OQ3fnmvblvKhVheiYj5UpJUeVEnxBijW0ZK8wlkNROjO7rIIZHGRxgCSE7NqkAiUYYSVAjsrd2b2J1Zi2gAMA1sWNZ8lvgTHH8oVLRrUOorXmnlIB+Za+Z8I1jehTpm45nEIEY/7ni2dJHvHJRXWwo/THnFgUWuEyW6XZ0AuYNXRxahy3XJrn10S+OUvIydDMZe1JyM2HimdCsSS45CInI9SknzI3df0G/ECSU78KgKOpatqjgHwcVxKN0e+SGbh66q6aRMT/WwIi1cJtnowUBOp+HmozSKzTr+GxGMhJztRUd3AuaESCFaeBLlEor578BEaKu1KAgjBTFcyd98HuaXLyG5m48aHL2IpMHFxrI6giGKLNfTRCvlmJEFpyjLAqOhlqz67YpWDk0IHXI0XP1mrXRnCXOmZUa3KBBLyO4LBGu40YllvEiz8HSTKqnMQR1WcLm1PF/RmfCbo7c4WId2sr9V3p7uqBFVo54zsJnNQ07hle7o6AYy4UiKCOOBLoc7OnK6watxjIhEb0Xecp1Pg9yMbRUA9lvlRLz5i5eAITp+Gh64cSLPSVNlR6fR7RQy5mPLvKxG4KZHYFr9GGwzEnD4Qt/XEhzdequzaehzub4Sa2wG5Qy6nT1H3hUiHg9QGM1jRhJldFFVJsKrCHlfRvoJTuBEaadqcIgkalXYiDIYbgqjnlCTTMoViz0jiMfjzwV+KmTmK8uyqs1LeT6flJfcM8wJELIaBJE6UFl5UToYJgdKKwFljHbALgDfQgyNAE6gmodyVHE9KyJsfds5SHtG5Huj242BVEAMwV6iTBR0TV6r7s6JJVILG5udcka3Vzp+Xigqic/RXqw9g+7EIWigcCeIizEGqW95Q4pCtaAFc9o+14ej25AHVJ5ay1I9L5UnADI9tYAiZ5caBhM0EWNEUch7bKTv43TyhvqM3CtIAHZ1PZGz+gOxvxzNmc9jfmhdEIretJBfClIVB5WfjC6rgka32GmyowqIrGeCACn4iNfJC3mJAgdlCd4AACAASURBVBMWoIbLn1naZ1FCT2YSGKze0OXx4kRcITAKE7yaCaGlCMFeJpOM1B/8kqKGP6FJe0IUxorDsdcyqhC0jgNlKFhJE4lWrDQhc2ekoCAww0VLnIKleyPT74zd0R1RU34nv8AbfWINcliuzMUKnzKOp1sKYjGPhGCH5JUvOo7LfDO6rXPXalTmNGfQXedQZOyUbgidPgyBt1aDu20jorVxwt6gRplxyDzIzUV7GODO1lSL9f0SfhZReaGpMwi+SFtPty86/3K6k5OMdXsvJFCQBCWXJqseQ5b85R5bLEiys2VwDa5EkH0xJisXJLOAbKs7ZquuTSAQVYjUB2qksiWaYJNU7+6r8V5JYibsRL7LR2VSwRQ0ymYz8ZpR4pCPQNHVSKJ6u/rGGOk6VE9IgYs7ch+pc2NiDXEwGrAo5YTopiPPmEG3GCEI8tb49JchID2ZCObRffVfopI+B7CGMX+NpiFcZYcYpnsBkDr4nG7xATZ+3eGuzombvKPO0cEP2PZnk7agc5Oh0J2f3CW5dijc+1g83WRGLUFJUhJBTolfgkR08vbj5CPvsxVa0xB+9U9ucqhWdEnlC3NA+gIscQj+uck2pGHPDuXlt+jFmjlrcZoOvcnKShZ4YejceBLVIaSf0v1tMrJgzUhBvvVIXUEO0w1b9RPZxuj6TskPGq2ZJUMPvpBjOlLXaWmRkWCuQvsdBPJGP6aAS9LnynMCn0AlDA2u0puoT3fJ5wTgnFWr8NHfuA333XMrPnLPrVg4u5P1yXtSR3fJZ0Y0tuDW9VeYc/TfS3EJQPeCxbh29dmwZhfXARvF6Qj9tgdBeHnbLdeh8AKS30TKp8DblYnnYadjmQyIEZIokzgkOZVr9qJluObi5RZJpLjI/9OuWnlXh9Lt6wfuBKfo5WMyV7rJRz5ydKfnNja3Y9XKJcpXvee0dIOjnNWDVEfIaYrwX3VGxmnA7Tdf5WQi9zsEUEe36rWCGIKc2fLeG69De0WeVSdvV4TP/i0t3ipfpOAWoYFB+BT4hH3i+0mfLzbFu8PJ2Qc53XcngZmuiR8Ve0m0W++I2anRbDqc7hV6Sd6Oa0tAsjwDIpQxdVmm79hTRtenr5C6ZkYoCuScC6jUdMPeU8mx3O2+04NlNBpX2FhrbAik13pxCqWiVEuWLcOLGzfgzcPDaGnvxP333IB//uLDjhMOuWjUKhGKCubP6croBhthyfsIEEs0Nregt6vVomWENeSIsLhybktnVo2ev2AuQiCU+sYtZA0xgSoclTjK6px93u9ZQU6GcvJSiRPHDmFLny8WQ+eclJcVh49TK2NVjdjefSx1pchRKiJ763rmMIRuO0HL3ngf0djagdWrluP1tw/pnH3/TFoetHEjokM/8jOj8MZH+adUI/2bUMYpPPnMi4pIrJgYcvQJq8Foca+uNgEQnv3Fc5isMV1Ejm7BpBy5S7MfW8olVTlDSBLZAy/QOQN29HuqjedsK7zqpcVIpLlH8Nvm5V5Pn9wfa+6zYHQ755xMtqZjVLQgVm+AWfHI1lyT/khUd2vOSNBYII4uf9U3jLhlqfplI684Co/k8+wUIWFDUO9Ynz/XalXUajVMTk5hYnIKlYYW3HrTWgREzO5uw9f/83G09c7DPbetw+jYBBoxha9/dyM6Z8/FvffcjnkL5uK5p36Gza8dwB133IBGlGhubcFLz2/CAMTnA5deeSUuPX8JqiVh35uv48lNb+AP//BeDJ84hSd//CTeGRgFALz/rtsxp62C4ZFRdLU2AiBcc901WNjdAioacHjvbmx46Q3c8f7bMLe9AROTk+ic1YovPPAofud378XIqSE8/eTPcclVaxDKabS0tuK5ZzZgX98o7n7/DahOTqK9rRk//cnPcHhwDIEC5i5ZjiuWNGO4eS66iim0zerE0jNm4x//+UGMTiWDaGprx2/+xq2YHJ9AR1sjvvb1x7DiotW49NwzMB0JB3btxBPPvYHf+937cOrECcybPw/bX3oFcxcswOIli/Hjx76HqVmLcO0F8zA6Tejp6cQTj/8EI01zceHsEj96bidaO+firhvOx55+wnnnr8S7du7DRNGOyy9YisnpEtWxIXz3iU345P0fwujoGF7etAk79x5FoIAr167BkjntAFVw7OA+bHhlH377/jsxdGIIvXPnYseW5/CzF97CB++5A51NARMTE5jV2ogvfO0nuO+D78UPn9+NX7t8GSbLCs5YtAAPfePbODA4ibvvXI+piXG0t7fhhz94AqOxGXfdtg5jo2Noa2nAY4/9FOtuuRFN05MYOdWPWUuW4yffegTv+427MTY+gc6ODkyfOoqvfOfnuOb6a7Fq2WwMj02iq7cL3/ji1zA4ndLKtImMlzfZ2UohUVMNRdlib17PfQ3GCsAaOKMss6fv9R23cOhZTF/TcIf4BW/Fml7nUyRLsYGK7XFPEwpFhQ25bqWC2Dg5EvmIrnTJspm+7QmKEjRtQPKi2eGrsDV0dR48aVl3z78XUxVkYMtG8nPDTeuxemQK3bPnYPf2F1GrTuLJn2/CvNldWLTiHLxr+TxcfM178OB/fAvjUzV0dnUihgraGgO+9fAPQU3t+O17rsXJymyMHzuAH730FkKo4CMfugXf/8VrAAU0tnXh8vPm4fNf/jZAAR/92IfQu303Olsr+NznHkPJcHDhWeegZeI4/v3h5xEqDfjjT38UHb0LcFZvBd/6wS8QYw133307VowQ2quD+OJXn0NRacT/8Qf3gkJAZ1sDPv/5R3HRmqtxfPfr2LTzUJrLPTfh7WOjeG3LZuw6fAqhoQkfvvM9ePCbP9ToRQRQ0YCTx/bikcd/jrXrb8TKJb3YursfIMJtd9yIH333cRwcHEVbeztCYzuuOG8+Pv/gIwAF3PuRezB7+17M7WnDF77wVVRae/Hnf3gH/vJvH0Rrz3zc894LsGn3MI4c2IfvPbMDoaEJn/7E+/HwU6/CzjZJctz26k6c2VPi1beP4nc/dgce+OpjiBG44tprccHSXnR1teNrX30Y49Pp6LzmWT04d0Ervv7dpwEAH7j7dnTuPIA5Xa349y/9J2LRhE/dexP2jTah2r8fDzy9DaAC/+en7+OgnQytUpvEl779I8xbuhLr3rUCK5vm4aVnn8e+40OoNLbgnluvxSi14Mkf/xQDI5No656LW29cg9FKM3ZvfxGvvH0Mv/7RswEA8+bNwf/8/AMYGpvG7/32b6ClvQsXLpmFzz/4MADC7/zB/arzkfLVvXz1DfqdYhNGYWXNXl2JCA2EWoDXVyjweGprgkJd/wyllCftlOVl5eiQlqIZmZuZErETK9lpVch7KaWjdGcIMjH8OShtpClLXxiTPgkbR9MOkMK2KGtBho/s+rKmqAQCLQHIRjHdFFRfufbHxjuhPPmTp/DmkRGACB/7zXtwzsA0Vp+zEJu3vY05PV3o729EEWuYnE4RdujUMBpbZ+HI0b4UAaanUVJAb28Xli+Yi8qsOSAAB/btT7snEdHa0YmhwQH17McGRtAzqwn9xwe5HkigQOiZ3YNjR49rSjVwYhgdXZ1YvGgh3nPNJSAinOg7iq6eLhw9fCyJoTaNE6dGgLLEwMAgIoDZvT1YsqQd7XMXA4jYu3sf5iw7BwuaL8SSlVXEWGLXrt0sP3dKNUUcPNQHAjA+PoGGSkWVsae9EX2nxhCIMD42hvbehRga7E8KV9ZwbHAEs2e14Nix44gIKKfGceBQPyIItelpgHfRDg+PpXlXpzBdk1w6GWzQk6a5ZlI04YyF83D9ustZx8axd2waQydOYGK6qsGlo7MLSxafgeuvvRwEwqnjfYhEOHKkD2UZAZSogdDb043Dh9/i/LuGE6dGISkHATh46CgIhMnxcRSVXszp7Ub7xauwfCpB8Td37cO7r16Lyy57N6YjEMsSu/YcxqLze9F3/JTVHULA0IkBjEyUIERMVWtobZ+FkwP9queDg3y9D17kdF0LypbmBC1sRzZqcyrR6byccKX7RnRMsKyBWEZQEVDWfLMddE5WXHfNiXxdKjpX1EGJ1wgUUIOcJqpEpX/aYTeco3lkoJ6Gs8fo/hOYJCmKQygl76IUj2hNXnBjpE7HWJYp+4ypRbgsa+wHXJ7qimnZ6gz/3djUhJaWZnTMmoXezlZ09c7GscOHcehoP0KlghACdh8dwrpLz0Fbeztuv+29aGuyMxAl7dqx9VUUDY3YsHELtr6xHyPDI6iVJVrbWjF+sg8dC87EormdmD1vHi5Y1I59x0bYZwttJd7euRMXX3kF5nR3YNGSJTjzjB70HdiLU5Mltmx+Cc9u2YHq1AS2b9uBd11+Gbo7WjD/jEVYtrDHkCOAl1/aisbGRvx8w2a8tucohk6dwuYt29BQRPzsmU3YffgETp44yXKUjlZNgrWTUnNqAM++/DY+cPMatLQ049rr1qKThtEx/0wsnteNuQsWYtWSWdjbN6LRyO9pKN0KzGWXXYzuWa1Ycd75qI2dxOBAP1asXIHWlha857rLUESgLEu0traivbGKnfv68Obrr+PpDS+CCDhy/JTyS+Tef/gg+keqeOmFbdj4wmsopycxPMHNe2SM2bnjday59hp0trdi8ZlnYfG8WclIeKWk/lSq57a8isZQw9O/eAH7+4Yw2N+P57bsQJwawVM/34SB0Sr6jvWZTgvdMa0KJISb+Heq7xB6Fy/HGXM60d3Ti/PPXmR6mAhSnpUln6QdSwAlnygeuW5ScwYq9ZOQ1/R0pUYCLhmqJlv+ltpV0PogVB/k+sj7u7I9MLrCJrZntkBEVCw/56I/C0VDgxZrokB77x3ZWfiUgsid5Ufq2QT6gdjbEcHv4hNoRbDzHq0HIH0dAr9fRCKSe6cDUToNG2THmRFsaTJQAQTg4osuwMoVy7Bi2UI8+dOfY+ebe7B4xUqcc+YZ2LZtB4gIz216GXMWLcOlF52NndtfxZHBYRAijh4bBBARCNi7dy/2HxvG2isvRmczYfPLb2BsZBhLlq9AdfQkNmx5DVdcsRpnLuzBd7//M4xN1RACcOTogPKhNjWON/f1Yd3Vl6CZpvHSzoMY7u/D1jcO4qo1l2DJ/G48v2UrJsYn8PbBAay7+hI0YhJNbbOwbfsbABEOH+3H5NgoDg2MYe2VF6O1qOHFbW/h5OAAhqYrWHPZhaCpUWzbuR/+HSbVyTEMDo3j5OAgxiarCIEwcmoII+NTQIzoP3oY040dWHv5hTh+6ADe2HMYO3buwRVXXIKl87vx2PefxNjkNIqiwOEjfYkvRcDRY4NskCWqRQvGB49i8YqVmNNRwaOPb8D46DCmK2249MIVeHHzC5gsA/bvP4jueQsxd1YTfvzU87jwolU4b8VibNv6KobHqwhEOHxswPSprOH1tw5gzZWrseyM2dj0wnZMTtVAFHHk6CDrArB//0HsO3IS1669BOX4KbR19uClra8hBMKRYwOYGh/F4NB4MsLqFN7YuQujsRFrLr0AtdGT2L7rII4ePoSivRuXv/t8nOo7jF0HjiXE1z+IyWpKC/r7+lGCcOTYcQBpjkeOHMVruw5izVWXYk5HI6qhgp3bX8NUtBUSXanjbkxB0DPe35HZkZz/IashbmVFdzSTjiNGZXYVpeSh92mfDODqIFD0rl9GayQUeyzLapVuuvPjo5WGllbrtYCLHuIrPBwyjylPsIq3eEA+D4CXsqTgotBKUhSi0/6t+V19zcP1Y9hkPeLQOArlnHpGy+NSnYbfmsX35xV32HWaF5IbS+guNHolnkcV4OnploIVk6ArUImgxtYOfODX1mLr1p3omb8Ai7sb8O0fbHB0K8F6r84VrmmHoJHQN+9I7aCse6+pbyISNJhgdXCf1TTdkiKaFL7PefelWEADeOaV/Y5Ovk9RH5kokdMtBpHvvAW0WapOH7P9QgBaZ3Xj9vdegle278K8MxZjdtM0Hv3pFhBSNE/is45Ve4RDo6BMtk4LoGlDsEK8pgxFIz5w53q8uXMXKi3tuPS8RXjgGz9U9H063YbSHZDptyp0mEGz1BUkOclWBn3awHapXbEE7fWYQbdc+0vpDirvqcmRcXUW6lq02moKLYRY85LIXzq/TIDZBh2vbKU1xvg1/Jz5UQ3Jr8OLwvlmFt0kJPcFMVBLbSxPE5ooY7ScueG9j6dbrs2WkrzsxIkguuYbcV7sXKSWk7U7G39kS7AsqbW2dWDFmWdgdOgU9h08xn2lvIzolEDo1lzVpX222U5m+Uvo1ufil8jbXgcYnV6Y80xzb+/sQiOmcGJ4wlRNa1r1dKdl+Bhr8hT4Ziu/ZOiX++x2V/hG1GjZ1t6BFWctxsmBfhw43K9SsmVKW0nIAp3S7WtwrMvKDyfTusBCIDQ0NeHs5UtQnRjD2/sOoVabGXhkDO1Mdc5ZZGBjOl1zc46wgr/wMkI2IJoDEpllQcoFmJnytvnBf07Gj+rU6BjdfOfHxypNbS0WoXkNl0hbbNXreEbHaEzzzoUflBmyTCKbrE9xuL9DCdSBXH+CCdN7R3lONne4iKRTn3n6sUW83IjV4XmEg2iKUicYHdN50uh4YPxx0V8iYxZV6ujOol8uXJuz47yjKev7l1UqH30gRuGfamgkG4+kvf5X0C0jOBSXIz4vb8B3NnrabUu7o/s0Cm2ypowm4wnzUeReJ2/voH413TXlZ+6EYzZPL++ZUVr4EHW3cP3cCHX38GNm0K4Bw9oGwL9CsOCTo7/S6I5REZKptbNv/inLmjo0ooDpqdHxihEmjVPc5FE6ZgMMTfkhopuOaWX026AZwmgmULeJiNMaM8bolMQcgETnhIgLG1vfMCVCUqq5lZivk1qJoARxKLoUxYWc6J7Jj5UCWemVP9q9kHtdxBdYRBRwxZrLsWLxbFQqFdSqVUREPPnUs1i6aC5e2Pa2KuSVV74bL27eihoBPfMWYmE7sOPtw1hy1nJMDR5GY89CTJ84giODo3j3JRdj35u7cNWaC/H4E5tMtgrjpY2bkLZkswxDQHN7Fz5421rUakn5T/Ufww+eesF006VcSpdAc+8HAY3m6YwPp+zqKEszDuZ/GSNCYQU3KmR/SqqvSCszK5bJHhFUVHDtmnfhmWdfdqgj8TnRXbN7xHJIKv7IfmQfidAhshceRKSmLlNV1i/iw3Y0Wnu6BTk7JM16jpjmDxmnsFYA+ODhHUzkZVdQ1pSmaJlrFj69SNxmGwiGNHK6OYDL0QFkqzDKN8UkFsTKMq1QBdlxaDDLFWRczkjym1xbab0zLK1dNcYyNW+RFCbBzLFCZTJIloq8DoCr4RDjFqfA8FuLO5DiD1/Ds7I3WTNdDpCJQgDS6pu+DzKejOmiddoJHXkpWby7iQDMfLlfFOTFzS/iPx/5MSbQiCd++AS+/cgTODVV4IKVy4RZAIBVF6xE4HFODQxg3bVXgogwMHgK16y5CNdcsQqDQ+MIRSPWXXYuhsYm8PON2zL5JLpltYkV1NMdIxpb2lAdOo5vPfwj/OcjP8YPn35ReUfk5O+MEdGK0FxaS3yI9XRDEVcq2glvTJfk3Eq5FxE45+wzEVjerW0dWH3x+Zjf26H6llrYC1x3w/UYHUivNjj3vHPxnrWXorOtCQSgo7MLH/rgbbjr1nVoaQgz6FZvIYbG48qhz/UggCD8gOmgfB5ZbnEm3QXvtlXUJrrk9zWVSb8TsChNp5Wn1h5QuBeM21mxri1d+WhNjyJBvQbSrCh0JznYlgkYf4TfIjuxDqfr6b0hsqmLtyCbg2dGecTAUTfxLU00rVxU9HuAuBWVnxvAxT/bIq3QlABE9qAK6Xz3KOALPsISjTAiWbVh973CSfaeahTgv/MGMoOnZHOKbk48b/H0gdIqjaEb0hbckpFYWaaoWi1rKMg5OI5I+sZqEGrTkzhwYhpLZrfhwEA/mubcgPLkO5gugeWrVmHX9q2gSjM+9IHr8JVvP4X337kecXoKra0teOZnz6Br2flYtbAZ1NiOpYvn4Yv//lUcH5ow5AH238y9roXL8JFbVuPk6AQe/8mzWHf1JYhEaG8kfPPRp3D9+vegraFEpaERz/1iA65efz1GToxg3rxeNJVj2H18AosXzEYc7cdXHn0ev3Xvejzw1cdBocAnPvI+PPjNH+JDd92IkaERFJjG9360Me2hpUbcd98duPDsBfirv/ocGnrm4CPvW4dnnn0F77nxBrzx0iZs3XUYFAids+fhrC7gwZ8ewjkXXoj5LSUOHR/G73z8A/iHL3wH991zI771zcfQ3D0P9951Ax741k9Y3hb5tZ4FIB0k43XD0IGvkUgRXBsBQaAimB2pczF7IyJ+N4nputdZQVP6fGkNV2RtOiptCxQMrZL0V0i6J2fW8hiRHbTqcRDkVWZ0K2+IkL2WANBxS6mLxPSG+FqVUrt3Yqicv8AvvxXsiWhFtQxREBernSd3OZ9tw5XGLCskpmdGmQsUQs3I93KY5g1VPLDmyGUV0UkxyPZtQhrDtZNEYT5gdJdVQOYVE2xLDi4xUCMsUTI4d8Kz5o+QIBI18ggQMedn49hWbqaVCL/Y8CJuv2o1vvH9jShjTClMjFi7egW+9bWHAGoBEeHytVdh76tbsWNvH6jShN9433V4ec8gqqPDePixZ7DyokvwrnOW4OmX9ujYqy66EB9u6wVAeHHzC+gvC5STI/jat58CEPH0sy+ju6MFq6+4DGd0tWLFsvl46Nvfw4mhUcQINDTPwt7Xn8OPnzyJT/3e/Xj7yYfws6dG8Mn770GDQygRKYC098xBG03i0ac2YmLaemViOYmvfvUR/ObH7gZixJo1l+K7Dz+Gd05M4bU3D+JjH1qPbW8dRYzAXbetw0PfeASIEbt2vIY3Y4neeQswOjqO3oWLcWzPLpwYHgeN7AeaL0dTpcBUzQKeN4Bs9agsNT0Q49NAGEuVd0FBzySJkGvEQMHOxdXiKOiqmCYIvv4h/RC6jUGQD8xhlYYWxPg1oqn+80qF2FUIvEeGbVMRIoGoonqceGHnVvhtEp7u4GyZ/xcrZVnlo8qI3/xkuaoiA0QTtBi/KxbW7+nwG8uyFQWpeAcunqpwojGNvZ24oOjGEK9bCtzWjtBojkqQALsOrZg7RRHnoBCTt92TpEAkhEdEfvO4ujZxaN6xqaNwm65UWxk5BKA6OYGmtlbuO0nLaY0hoAooihkZ7EOl82r09PRievAAGjpmo3v2PFSHjmO8FlFUEu2zezrR2X0e5iw5EwCwe/degDpx8PBRxFhibHwClW47ii/GiB3bXsW3Hn9eHXfXwhb0HT+BGEtcuHo1FncAr+89gp7eLlQK4BsP/RiXrb4IC+fPxqYNGxHjFPc3FBgeOon+E6NAjJicqiKQOVbZhTzcdwhPbG7A+vXr0DOrCQ995wmMT9UEbCbuBMLxgVNYunghDp3cj1k93ZjfOwsxlrjy2nV44+UXcGo8vVI9FAG3/tp6VKrj+I9vPo7WuUutpRxJH8pYg3Y5Or0RHVe9BsBvOVZ5e6etY0ICt52jKkhcNY0LyLLnCSGhEj2s2CHUZMueA053ItL5thIY/ZzVhkgdWgqg3OiodTmhm50Dn4ciWw8UUfHfer9ENkc3e8NU+yPwu07ZgDykEkZLtNB6QRYhrfACjiziMaWxShpL4PIm703ls+RL2AjlOma0NK8EPnSlCBWXe6U8K9TlZfryJBBCUeGt7jaGXV/XuwHxxtb4YjUWEXwJRUOOb5oTSpOZSzsIAKqTeOdEFVdffDbaWpqx5ppr0Hdwjzkfltnm7Xvx+/ffgc2bt+OF1w/iD++/HRs2voiCX0BDRHjppVfRUAF+sfFFvH1wAKdOnNJt7LLNW5vbkOZVqVTQ0tKMluYmtDQ1QRI2QsSCBXOxd88+HDt+EpVKAxoam7B88Rxs3LgFG1/ZjfNXLFLHna2qaE5fRdus2ejqaMVFqy/Gwt5W9Mydh4bqGH7y0w0YqjWiu7WReR/Q2NiASqWC5qZGbN28Gb1nnot73n8jrll9Nt45OohZvXNx4aJ2PL99HwqW3zXvvQ5H33odTzzzIhAqOHHkAOYsPRuL5vVg+Tnnohw9iWrJ8lbEbNvW4WQhZiGGRV5WWqcxPZRAEShYYZH4ZUJyRAOPKkdR+p9M17IvRM8L+K5LIkp1ENE/adoSZ0Cm/+k9vyHxidFxVhdUdMB0O8elNSUKdrqd/p84sQiiQMXK81b/WSgqDfqWdGekSghx0crDJiECpMeQ6QEvUTanIXMUkjKkmfD5FNmbooJB2bpqrj80x5ZJYc+ACFpkK7QIanHekllilfA6uplZSreqQa5UgYxuFYA6X1FWwvGjfaim8wnx1ptvY/6SZbj83edhuP8InnpuBzt5jhgEDPb3o6CIV3cdwMmBEygCsP3Nd5TnQA1vv7UHA2MRay5bhYY4iVde24OIgNFTJzE0lt6ZMTUxhoFTY8rDs1eehbOXL8XKFUuxZEEP3tpzCLXqFPoGh3HwwCG8690XYfH8Hry8dSdibRrTRTMuu/h8dDSW+NlzryIS4fixfpRUIBChr68ftTIhxb6+fhw4dhLrrrwY/YcPYvfRkzi09yDOOnclLjxvOd55exfefue4OverrlmDlhCx9MxFOHKkH2MnjmPD5u0Yp1Y0VYeApja89MJWTExbU1VvTyeWL1+GlSuW4qxlC7B79wG89uZ+rLnqUnQ1Ad9/4nnUuL9D1d7pkV9ih4Br2UQJaOer6ZTTLcn/JXpHCxTeUYiK2QE5ojOi2+4IB7YjUTh7lju7QtC4Q8ZyxqYaPiFPXaAkmf7LM1nPtFNUayH5sq8UgCXwlbXpafq1998/2tDc0Zqe65pNFO4kgsuyxg9IxhVCBWVZ1QcwUFK4F0KRnexjGY2LxhDIZfURE2pIYymacV2kWc+FO7HJp0OOiVnOJ9e61MXTHfQzl8uqICMoVFDWpjWyytiebls6xP+GQC+POwAAD41JREFUbmQRyNMtwpRx5CBdcdh++VfqL8pHItjLnMW5i0OTpeCoPAVg847GD8/XpDBVR3cau2T+SmfozL4G0SdXq1EHzvWBogF33nkj2hoIsTqJh777lL4wyRCMLNvH09ANfVamD8JnpUcOI5ZvU0CQ+dgqnLQ6pzlLkTOxgnlXlgCj21JqTzxmybm/9TRA5R3reEQAn48qL2T2I7E+SHTX4xANGwkqtpoL0x2Id68G5YGYmGQJeoxEreYCUdQ2hejork1PjNNtd31yrNLY1uLXcuvX3G1Diu9eM2GL57QCjtikjOG2nnNUti60hDK0JlKPKMicQjocxRkXoluelflFjfw+B/WNVqq0roAZnQGKkwiy8UryUqcScm2qf4hQdNbKS1M6U1w/n/pWdL1ei2IlQqUBsazl18acbvu30e0VyhuQdsoy3Rp5onUJKg2l72GwpquMbsfXjG55LaTQm+ClPl/m8r+j2/NcaMjlHWbyts6peV21Sn893RXTLFklc3TLfgk5/HimrNOYvp/EYmB9T0cd3co7r+e/mm7r3hW94HNZCS5ISyGdHYY6lcAvabI0W96YrnTJtRQwPTk2XvHVXBABZc11TQI+OlEIoBhUmCBKR63JvnzyxJvTsdZc9uAeUSgmkTnARYn6yBQzh0qANl4Zw9MXikrqYZyLeMkfMmoQujkyU8znX0qhUyMDZQ0z/sfuyw/RBUSpoymiGI58Hk2pE89J0QcFcVYubRIkVE+3h8USidSISSOV0C1LhdZ+noxHTnf3DUCiiGkedXS7NNFQU2C2cyEQoiesc9F2Y4oOeLr1IWpsBuMJEaCY0Fhhy/deN8RiFWLrMr3wQZZIJTUOKH1QkzoAvCNWqp0jgRmkRz5c0CTY53YvFHkn/tZtPyBLlwVRseZogDO6KXPcpHSL7cgcEm+LUGHHyTZZFLyiIg6KTI8IqCDGqJPVwkdSSjm+X1GHQFtpLAE7CB+VhVEsMUEcyQad8MheKJP1Msix+a7OYCjHORePcqXwBvGyUsiiDEol2mR/iUUCFYxEkZINyb3kh0T5JR0haAu0Txm8EeeH9fDcAilE9d2nUoSTTjuTuXO8bCQqwLpUQiFmFo0AROEXG1KMFvIyRCAOQXjJrc4OOnsU5LdAS8STVLRebsmJyBbodK06ce9xeBR1npC5erpTD0tGgvBY9iDxfTZfq2dZ7SxxL2/R5n/Lc8h0KqObdThDClFea+hocfJwknK8kROqpBiJTHaZW3LISXSJmI853aTXpWeZrmddm2Ryk7TK+MvqRRB0FyvIijN+aq4qnCl70L7xLMdSr+bqAIIUnMeTYlBqITWE4fdzWFStABqNCHKWpzyHxJjFc5BsX5c5JedgnqUORTmH5KSo6EW8eoQcPGIePY1hgrEIaemORzMSZcooBbs6ugHOI6O262pdA2DFCEqbtpkrvxwsJkMcFkDr6CanusIngb3MPnPwzJNMPazSbnQ7J0dyqLAYNTsadbbm7WWZ0Zb9nAMD6p4DXsLkRiNyz+SxhF6tJ7ham4swaWTmefbGNkh0ZROW1yEqmhEdMcendTspbHujdg7R6OaiKacTMaM77RTW9DUY6zXtUnGxvDn1iZwipUBf3/btgq0uLASjw8UggukoElKlCmYUhMSzpahnxTC+uazpaMaDoMogD/YC95VcYpeVxkqNUGqIJNBKxmUiyhormRHhI6o6D2cMupojqIUZ7ZXG4CArhENFzv9AIoAIRx6jkSBdwe+AtTlFQFO0QGSFsLIGhCI7D0QhpYtgUjzUKrmLOvocIkVjxuPg6HaoxMFdk5CvWwT1s/qH0C3PIgkirqmM+Sdz9GdJqs4A/IIn99pEZrI0AwmSKTUdId4+4IuUIn85GMZkqugnSSNDhCnF9I6U61AlXNpW2ust5TUV/FNwV2M+9yR34xupX7XQHDloWzcllO/pVCxFcLANX3JqvewQJtFdOS+GmaHyVLTh+izKWnIimo7YqyB9DSZG0xnfpAVEFJyihRBiBSDKnIFaCE/AKaBdBzEPU1wPx/i3LvFIOzkRR4OIWHMFJYG+lA4zEWcjxdWIBLP8O1Y1ZfFY1BGr8zjNeaDeQI3XQjdX3WfQfbouUDUV3nrM0JfhnFW4Q3KKSB2yVkiDGkVQpJGUVrdxixHDHEUqgMWZdIvwS6u35EYphuW79hgVykqBM3QDSQYrsnqKr9SLYwBARUV3a4ICG4TslDQvbEVhzaQVZQgykDTB6Habpzj9FP3TlDaQ25jGzValoEpPd7DYIc6O5+IsHoAURc1IJe3Q4qDSXUokRrYVQIKYFPnVVQOktSx5fWCqLYjepZO6bfHA0FGJSCG9KZ3TkiiHaYvE3M5xDZsiK4Ppoo0aCOQ618xG6S3q7gUlRJbfRsgGKrfsJYYjhsET0CgZUo0iOA+nMBIxoQkA1vPuvKRiK/nPAhyCrVMnBamIKsAwmRdwzJZNk+OsZ05U5msBiR2FbNoRur2MsloDCyGAVGAyby+2jG7hidAN/yPIhu8mLxMCsaMQNGWYUWQSoS+kJnuhj/GYjQfmWC0ig/c/RDc3kbkZjgglJUYCv0n1wNOS0CPBv1RZHUVGtuTMVui2Va1oAUfrQ241Lab7tV6FiCJIXUjQCBzdJm+/IqDB4JfRjURH4LeKRUGzMMeW/ik1OlmZgI1L5PTC0206kV5ETOnA3FCkbmNXQBUWxxl0Q4u1ku5oIOQb/JGZCZWGHBTAipt+zkBEhUAIRYNbKuJb1HjTpAyeiLfOK/I+P/NLhXKt/TD3HAKxB/OOUIcQkjAFInF0JTcOYH6CIafMyXeYKrRyKMYUwvOmgOyLyZYVNdLaOrc6T45mBFufN5q9kclcpSDLGsxr8bYk6k+NAnyFHXAIJDrH5QxcV1QieEWA4avku+R4IjIU1BahrfgS8WfQLTISDCjOw7U4q/MSrwni7f4ssEga2S21zczItfWnOcmtSUfkKjNkMRCD4+ycS6Hbp7himIWpkNINRDI0lETEz4ycLjhnJwFSHQqjSzE6X9i0WhTpsnTk9EyuT+fV8kQ1azFeeoQgaGXGUqw46FCkbQwwZ5RQj614lqWhxTSv6FCR2DyhEkKIIYSsSGiQ1Xt3UZ68AGU5NbJJq1KoceZLmOmQ0liXWkRI5TY9s6bQ03LFdHdibL6+rsYn8JvnZOCFDVYhsC0JikByui3HE8WLIKXDaIF+FkUg0sGndEs9R4p0XGdgOMszZBLSMqA/FUtI0/0CBFidCNATqQSya67q6bYWdlWQzGnzPAvbVp0ZihgkJUxhtS3jve9rkOepE4Qd0JImxCs/zunaKw093VGjospVImKdUw5yXoRDyiiEdpi8JZp69FgYzE/+v3BBxNCrTwHVxDzdfF4suLEswt5OD9WYXE/lR5GAonhxOKU6IaU7QvlUFOZsxNGHoiHRJfWWIHRHnQYR6SsCjLeFDuOL7QEAlbWqTiDli6URxOQCqUAllV5SxfOnIpEqYygqjAiEA54pIiAPo/lJriNQIJF3CGLEino4X4vOSKyVtb4wBo3IiFGX+GJZQyxL/rejm5VCOuEkquZNQDJ2+lzOIcjoVgcnkZgLwqJqMWawkIi4wGYFUOWJODY+wMTXMbyBaNMbz02MQOgmAGWtqjJXzyLXga9zfSwhSCHP+iskjZFzLORziNuMEgrrdUVkV7JSFjY2UEe3608RJ1ZKT4TQLQ1XNX3DmqWPETHWlCdlbVrlLvJWwCNzCs7o3Fv0fGAMoYC8XtPlFY6HUJ2xmhg7LP6n0OZ1TvTLluSjjpfT7ZCK71FR9J90WlCZ0A3nvHXWjO7SXi6oTNJEE30VzWD92q5MoCwB9vSAQbZarapQxjo/BSmw53NnXZTa6JVQSYI61Yw4IzYZWBmT4cux6z5/BfyLZ6M6gXSSkXWJiuePMe+eU+HEaJV3DxXLks8eYBrYa2v/veSFfmmKuAJfmpJHyPFmpmTW7WmK7OlOtBZqROaYapniSvph0dEKhlnFvRQlJTVk2TGpaSLruiA7eV2k74NJ1yae2JFtRmeqozAfyXpJkpOtcWQL0AKiRGZ1iD54cAGQnQfI9h8p3S4ts7qLoCFrCwcJ3b7/I2+mk/nIag1gxVJfZNW2ARlTC+EutRW6Q0CsVZ2+uYK61sO8Ptp16ScVuRNgiTZP1TcgK4x6ZyIOSGNEcorS++N5HtlByvKyvHYjP6Iv+YCKvIwmOW0ueAU2PnCxRTaT8IOKwlYx9ERrOKim4cWWZaw6Hp3Sx4yJyjA18ui8ukSLJDx99yjAuWaANFwFCubIyIo4Yl1pemZY6s2DguPk2RnKq2EUFaOvZFygAo6OPskQuZ/E9VLo/hqGxOQNwzmQ+nZiSYk83eIAI/zKERT9pPtsSVGUObAR6oqVoDvO7YuK1KDKTE65HIxuMq2EnO9o79awrkhx+lLXOF0z20x+EkdIOVIgAtFV7J2+EfPJOxl1PqSv8kkfBbLFLdaZUGl0BlJPd6oBZT0b+p0Zoh7PUDp7gA8GpuOGNJULblwuopZ8Pae0hrBI9SgFbk53i0od+wgobdUo9XRAl2IlTTEEXsycCzuPiiin1SXSRGK0rj2rKucRGIoqDFGoY/CQONY5FAeTjVG2jAaNVAIheVVFO8z8eH6py6KbOild2pNqNSnjhBZTQlvjzz2wKYU8336cE3O1B08XAF390Yio/DQUlHWbOtTjC8tUx1eZl5eNn4vRbZHX5i0ohDTt0Up6Tp7KJP/Jl6BBpmAyhOS8Gvlm6AJ0WVPkrCsU7ki6+rqY6Kv/LY7FeAv+DEjWC/suC1D4lXTrj+4kjf4CpdvXNYTutI/ELR3z5eJchCfpt6fbDU1w8vPyLxlJ2xiq3+q/UyCgUnjh6CEg77ZNDklo1GuT3cXKxPjw041l7XoKQcK8DmrsiJEQKKKMRIHcfv4oKUSMkZjZolrkC6Hi5d3yZGShuThAkRzhjAQIkNbztFwqKQCieEy/fIfIc4n8vWhNBM9RWM7t7AZvKPWc5D5VsBDFGEtipYwMDTzdaZQykoOZEgIgR5VRRiDfRemIWO4NIMi6abSWeyLeReiWutgtihJGROvrjtYwoXTLj3fuMIu379OkZW1C+AmikJ6cjD/xWN10BFGIIk+myzmgkJgD8nNWOSTxBQ56EWB5y/PSONZjcRq6meboDM3pHwSx5UvJOS+lrUouL0EUiEKIUi8xutU6CM5wJSDV0Z30R+ecuFDGkgi2Ri4F/EBFjLGkfI5RlEVkBqM76U1UeSKzPU0lPNoyehWE2PVlJKkZIlKMMU5MjD79/wH42csNqAsMrAAAAABJRU5ErkJggg=="}
,{"background-color":"linear-gradient(360deg, #606c88 0%, #3f4c6b 49%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/45-degree-fabric-dark.png" , "transition": 0, "items": [], "notes": "", "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nJS9S5L0yK405mDmNZn+BWmk2Z1puVqA9iWzLkKDgDscILPPVZ7zdVUxyQg43oF4MP6P//P/+r8///W//htAAEjcCVyB+tQvCWQCGQkAuPyrO5CR59q5GAhk3oi4kEg13Y1G/ZVAAnGdhzNvtRsRp0+AbWQAUU8EkBkRkeeejEBk1nM4zyaQ528UPRGZeZrAwJjIDETYF/Vr3v8Bd+DwDBERKHom+wrtwA0g4qqus74Fob3hBsknbucq2+JjGac9w43TcDRhdyYuqHmn9ae875LRFQAyKCtimLx9wx2SLXXDcft94uLGbXw+uAEUQ9hi5h8iPnF0Sridrmjepl0uDl5LhnnHud78O7ieeMdzdT0QgOg2PhSvCzeVsMR9xHZ0O6UH5HnpeXpXhz/Xv+AOUhdugwgA98BdAslARv79/b//z/fzX//7f8fnf/tfau8CgBuIS0qL9bx/DqrL/yrmkJ1+pxCde+Izrkcp0GnPlMVJGOQYPW1RQCmUhFmOCzSwvFtBB012bWN/+9BAP6QsTRS7jXjv1/iBf8XdhnVwH6ON4TF0B4C7+HBojEzQ0FAaiI/1XcpMxY0XWQMALiCujzl2OoRNcT97+q2HTX9j8PzZgiv3FWVyb7hJL507n4q6n3j5UzzHuHfwx75M8tHbyDfci1/C17YUV5rLLv2JaC+AlvXETeeI8tHTWWb+oR2v8ZZ0RCiWwNoYIfPC+EgPIvD5J/77ewwWLRcPMmB0Y3sxmR2MGfOZ2d5k/jGY8z8KllyQ4xkO0bXist9zZCJ9mT56C459Vd/XBRSDH90w6mUzy9uemPjg7K+jTuO2P/oxdv+vuMsQ4uDINOX0bhNI3JNPO1sL4mbTDMcxaOwsbVyoYONZBAYQRf26X3JI4AQhSFGHUwpniONm9zm/H+zO4knpVJhOJA7m7bztnizH+gv30VUpdLeT5eC9P2WKRr3R1I6CtL4EZcd981ni5nNoPSVNUotY7aT96bqr3KJyrInDZRMR+CqLKWFFfORhT5TvvqiwLepm4LnfmMqhjBs02hM29cdrc9gyFaUYRU8aaUIzZlBozpjVRwvFI4MJIT4DW1jzIUdmShvkBXEXThnUiryxaGYb5PH4kF7HU4riTnngrv7Eno17Onnn/XRQ9qjkEuWECrMp/unwesF9GordNpLh0ro1h+vy5v0D7y/clAmj9XVkUn1JgEMXA1kybD9UNsB2cY/7G3e1NwLHlrVjz8mP4SCdPwJrvEE7HL+NGBXQyg63E9q4L/JuykHD4kAHlLik49fJ1mUVHQ1pFMuDd2RZ0LK98xnn1z/9nfb9jEiKaPnXipD36jtm+91xMaMzh8nR1aelfjOa4V+wJZC3+WFnx23Xsmgj1lx8odYyGtx9XcrsvNmR9g0376shzM6ChsKUZsgpn8if+BeZEn8Drvstgg/c5Af/EZ8ZBf8efXoQeHEUsK/D+BOfwn3h0SezyG149XyKNu/f9XE6qkzHTfs4eLOM65FBvtjPyH4eH8Pg19jnQ4+vfgyUFYf/OzA0L0Ywk8rchys5ZUHc38Eso/HOGV0PQK8xUEHbKFSh2ONDvzZ+DyhbkBI7SEwl88jn7drFWWxDe1rxnYbqQmnl1ZPDo3/6WUU1KgqeuJT20lsvHigFfeETNu4NeOM+38+iXyD32Fu4C687rMTEPZzXs9+8q/ai6OO4L+NRk68MVhkAI/66d8hbF9e11gV3pWdYPIvMwwluPb//cLLIouf+M7kP0IXhN+4QPW2co6GNe3/kQH7gljwct+n4YMTCrWvl/IWbfLh/45YjTHyfVAeYXvfTAVyfckJh7bVSPYYX7mlG5Of3ue59+8Tke7DCD7tuXjBWVKg0eozndvsj6qyCbASqermwLO9uUWmk9IF2KNshBJ7394D2P+BexrNwa4joAWLjFsk2jSXcLsvB7OruDXfoOxaVm0eAinaDPxVw3FCGSIKQ3nEDU964kEPP/F5nBunNyZ7L/npkPYV7ZAWG+7rqEWZWxPoLNwPG1X2bs3/gpqxUW2EmB+Sq5c2a1Qo6pV9D3tfnx/2k54ME8EVcNb1o05dvnk+P72hVZMQFr3W0IReRD6cwS698HoHydIze9MYd+Ts6lIFXVG3xHwZQVmnDLNLd40qfvtyflwjhuGPhzn1vK6X+5hhaUeHq5+Rg/w23RRcvJhL99amocbWs2G7eJfhExLdwe20l7B+dgeHxbHDxnvcoq1Nmw2AzayfnObKlMbmDnMMfu2dkTWash6LJz+J1Ozg6M8dnxr+vJ2fo2Pdl/HTcdW0Uqu1v8goA0obC/Oj5N9wYjqJpDsTFWZxr8Z6sMtyeYQ95s/9UkN1BLnDllX8+1np67ia6BR9ufCXoQfBPZ9OKMpWxIiMd1R67D9oAjh/5PZV11AfuP3A8PpRd4/BTg5gMXLjH+NsM6Rfunx8Xird3N+7udOF22H4vx9xe92geuAEfCDfEZwCpGZGONrPf7TwcfmULG/cY6wIj4xxDwV+4re9hiHc5OtOLkVF0e0OPs9tOk3sHecO2ccc26Nb74BTwdqL/AXfef0uXzQ5y/RTN1bb47DrZeCdutw3Tczcr6eM9cAezDJvloZO7Thb4V866CZ0eljxgFCYt2f9MIO1U6GXJfAzm9++espp3dEVtlgNxtcN6pORse8+6NF3CNwp4v3B7VCLON6F6+47xAhVNawFUrBJjX3hieOsn08FBp9OmdRrWnnjGPqkcu5D3hnspcx6lmwpqPOaajk2HDzG8Dyswh+vHcKhQe+z3iNhT7/+AO01uwAtu/3DRWMv0kH3DHc7QUzOqR43qDffqT/cMXQ70sobqL4iVn42bJGf5F9dp1II60kKdmc6wp7oZdA7uCITWWfR4K4ywFuZggNIdB9weiNnBYwpHWAiC0Wk7EmBWbNqrH9/jdZNoMsd9xOKMtMLjZWmZUi684u7s4eCJMfNCehI9dLDipQc54SbvbApLCjUF33g4aWVpsG66wMWnc+rSeFSKHZFTiYYMk9w211HXaxgR+YKb96XTgKMDcorGH3+eiu18CM5iyJWUOlT7vDsu4A2362hm1dvcMbwbLjOluer4h57n6kfGCWBnFQu3aPSsoQLqI6yxHyP71IX4/Q6WfW9s3CNjb0ytY9uRAyzYZmZemX/mHdtThaK3Rxj+4PecrjtfHH9zUq1AK3pjyV9ygkevw2RPt07rWmGH8VU5nfaMo64ybuxhCle8KetRBlC4w9cIkJEh5nkEObg7DQytkXDcbpgpYxh0Kep7BIBwj4KX8dLivxH8MrThMAUTs/Aw9Yz1XFyI0o2TpvLbPLhzzZw5DZOogXs4LR+GpuFG16OmDvavswuLpOA6oUQHwqeeU//3su+h45vuiryxDPkI4146+GRNLyf4D7hHQd244HUstmcZZ2dHiZlxuv6azZijiPiYbUe1d8U34oo59qRC0TvWJEsmVGkmocUUrf66e2XgY7wlZiZ6EY8zePtUtMcFVPTsdlkAzfbqPudcXpqZCJtrjlxDQFCa2u2++bWD+w93lteN6PSO42e/WRXvG8iNmwKdmYxH+bz/Cvdf0dVyEZsUmrNxF4/bt9CRfVrZEej1I5CD6WnX0HOJQ0MO3OaE6PB8GGHDyt91HcNthnHwEreLqWcjGndnBcoiynuReuFmn4ar9aijvE+/M1OaS8oPre3w+m8Nv80Yj+Fl8/WBG9ZeIPOf+un0PhceHly3ZU/odp0v1v6BSVuKyS/LRDJvbaHIPBoF7lZRB0NJso1P3qankMIiVFffXekZveu54SisKPmqSPywL7Y35/D1WUWeHqPaEtyRXvmsCJOAu3GjcF/fQ/P1kfGH6CjcNnZVawHz6m+473fcIx00JXVl8bTWC7EeJV5wq2WrEWjpvUfXuM6YWRnnMYJ/xe01GY9mdOYub+UE5vwGgXhG9aWnjtsxgzpLxyYjwKIV7/J2XS/jHzOGzr8WUtuI6F64VTPAxARgrhQtO+loYI6U2ChrM3i0rOu35aBZjzm4w3gatbjN92U1liP/qzg6BaGbUApzGh8FraEQB9FzmetijCk0QU1r3/f6tS5wOWOaUTGf/THDkK4csZj5wB2GO4yxfd+Jb549vfFg4n6MXx13btwXchhXGpyXuswots6IovYVQdlNiCZFRcdNWiRzw62+Qrc9cTuesHteeBV9X2dTc1bop7wfY/KXKXF/VhX/OXsxckrd085hrAqt7Gaovgctw4Of9mH3AL9x6z7Kjrjrd2U7P4IQ79HQ6xLP0kYFkx5hzStP2DWQ3vZiGmAOIQCCehgCL9Gr/iGHs6Ei+zRsXY/p3exLo2kpymiTDIlJlwuX7Ty+w3qGuKcBa9qRQonCXRg8mvjswTvu/qnx89tnKDkVpjKCsRDoaTCTl1TCN5nd3YYyD+OPhls25NBNPUv0jps8WviUdcbku9O8Z0p+4fbh7hvu19+J2/oaX1twctxDd4jZ9HzUAN6c4i9Zv+GGtedD3jBeOC7Xre00LGjou12ralx9L+IbEaFKP7/wiLM6OT6GXtwjBRedUGDMNGwKCNC1vP+BiqvOKI2hY85YdANoQyHQEqgLIMsg5RvcWI3etwxkpJjG7IEbvWpvpbRMWUNRBZ0a3n9A/iFHfQWFOxbujhbPILymDtlXTuUc6y2EbTnE/BfciTYQtnv5ff18y7uLY8GM8HWWZmUdWri1Dd0+Q196dkv98pSGhbvH7tXnYwUxG1p88Szw8khrP6X/HggqqNzZiwIHbvLUMbzhTkjHSS9iLO7TkgYAI6vJnLi9zZHdmqxXYIR0+cpvZxb08NVhWqPuTX17s7IKpk/GCAF7EqAp1e0JF5FzdWGa109UhbHbuC64rFtg2+tCDpGG3qv+yDTSZzjdiQI4C2KK4WPeHsujm0G/4dYy344Gc9hD3Js2M3BXNtYmXrKmU2VfjmHgTqM9fuMpJe3ffzgbd6S+hmZ/dmbD5+Oa9PUD7byGo8qnbuWaNYirHmO71ufOGvZwTSxYAWbhbpQWrRXcNo4f7Y3gFouXTReHRI+VuC+4B+0Pfa57xzC1bRuZ8QUyuA15GHlktWdeKDbXXrwTL7tC9YXnGFIMQxvuiAi2LDh5axQ59Khp3Se6FnE/++GmmaxlvAnz/MV4oI1qZE9Ou1emLfo7HQP3PVrXx5Tdd/x1kepc863HcoTEnSisl3AN2gFoBWRlbqqzKMK4c3F5PzTc7g/w7DIDdBTz/iudvc04Yz4TVvVgwRx7BoD99f2Nux2JnsGiOeIcBCOD7LUdc4HT1nN3lC/4Bn32PIdiYFQ3ngn3+TuEezluw63DbTSsRjvVh0MAfCn5xv3LVxuzpnMzOSdqNuR5xsS5ec4zr0iVvpIRxmCLJOFtu2PBvLf9cIMaY2IyLmyfR7mJPIW20c+bfoNtchzIyvWk4Tdub8ajneMOsEj6wP0vZHXlfZLiuPteLpgibn7nCvcIhU/chXXQMOpFFtXYxs+aQrQTY1QcMwJY7QgZZLxgoHDcF1oslkVgyy0Md9rvpnOa2SHua/TzwO3B85Ep/8Lt98ysVrEmiPRlHYXomf1wnUlohsSwezY2FKyuXY7b+PWQN15wzxLANyJSB9eIXd3rc5OU82pFyAR6kxE9rBO/XdsUxliNVkOhtLFV7yCNGobE+3NkysPhDOLNFXiE27S8PfqCQT9vIOOJ208vWilg+tCu+Ni4E2lTbr6rcq6evIVr7ox8p/2B+5H5bYcTU3QP1+cneI0eJzazmo372HgPIfL+x3pzWZuBeb3lgZvWaatf+aTp9Z5ebFppWC99qpsfuEemjnYcaXLL4/K1NkO4Xcb/CbfLe8mEmZslA8OepZZml8IW/bPalesOEk+jV3p8WWZtKY1mR+ynERzyuisKeKGMQGJnNxYJ3dtv4xffjEnRtCm6lffvSGUrMct4maU0/ZbujzpNPHGLGMfsHpvF1sJCGsYUrNE/cBvfDlhFTl845NO+c2Wmr1Jc2Y7jPhZkuIFnUZIRCXhko+HrE/p6O9bCHQFohaDR8sOnD9x1/1zaTdy3/T5xe1/Mhndx24vhb7h7Ve+qOb1mqHTCFiDF/xjPkpaJ0XADpuc2VT7k7Ssyr5+4deqZ4x50ekamNEhtfQ9v1qwE00jOTNjaBC3gKSLnaUqJrtJTGQut1yNy9nHa+TMZmFHRayq1NeZX2+buJIDGwgylBcnn5qE4T9xjh6LS23zBDfj4dzsdNi9Dt+p13nf7WB8neqYQARmD0dIpbDSPLKtDnINqRrvRqyJPU4xMRWdNAXKLe+y1NaWwPZNVRgQs43uZMbHCnfghBpfBD9wcfzvu+wfuurfw5m2YZARd3Mt1ePARzV/nWqrtkGdzfc5v3DH7U8EQ0FSv+fjWbePVxh0WgL1/k/d9/yEicN/31Dn9loV7FvzlRFaOGU4bDm++mTfCD/3gTagijf7miLK8zUiL/HmyeKV2nn5ZHwP0GMLUPTTyURN5YTjbvpdRrbqHM+nxWbiVPWzcEfPMDf/ozyinktb2E/dcZwLMVPqFdvFlOUSPCJ6BeWR/xc17b7WtKLWPe4bhX8GlWyVuW7MhKM67WLTlC+5cP/mVGeIIAJh0bdmMe7J/Ltxy9F7jUudpv6YFIbKi+Bwud+Je1+B0LJ6S/mFehftegROQHsXA7ba6eKMAwaUNTU+kt89WA1+mLcfx/Q3mxPUVzZPxYXPi/K4cirIE846rIPg4+MQKXDKwsD4VbVxwVf0HRrT22YLzVY/RnitGfYjR1w/uXLg9kmFe4+O5Mc7MZeA2GuiQn9N+jpsKZrhH1LX5fXdq2JvWiJsyMQMd07j8fg+TFu7Fh4nbnSyjIYRxHnlghkjHpelwyzZ03wUED1vS4n054DMb8XS2z125G7ddfzge0x/eT92l3pMPYB3Q1jpo6ErdpCyz/w3cbqykwXHPfo46bAcfx3Ft3Fqh7HpgOj4+5/qZOqWT8AgtZiweAmAR79kgnoIfjgKWpvGxVqw+Hdwtav8e7Rw8ylmRZ4zlTUEey5eTztEYNtY4bIw+Vl7Rb/FjznsDY+HbwrT2YuL5+YEbUcOYjbvaYEr+yPJW9sUfwyhhbS2nMgx78mGfcdFrWPwZ8ijfccs/uzN2mXBDFJ0vF7QVDcS9C5dvuOt+OuyB24ucj2xn4mnDd2d+7tsLC2fAcN0znHrcbbADGKfZu0BZ19+Krca3x/Wh52/yPtcDiUtbuh/BxyLm4+PFvR2tjZBhWOZNBzO8KHXuHRunfMprOyFGseGBVzSw4t3+7onbGPdWw1H0fMPtdLEJMwUujT9aOdoYS+iFexfNXnDDsyVX5qVw6/c3d4Ti/dNBFj0AuNlotmnOhnRYJvQT9+Bz435O4088PPbxmSW+BKddu3r7HdXWWxYRLp9/w41xfweoJ24W2eM/4R420rjPI5euD6z61ZzPcHjA5BkMtzuJLcfzzReMa14Ie5t6e3inp8fUsyLCo+5rimKRvKKDosXKcLw9o20wObkJKDAXZPHRjnCc6/4f4x6Leu75nejn9mR+vaNvE9PRtqbeHpnKG27Ad4DKMeXz/ISH08jOX3TWAft8iy7jWhpufnfpd+Ee2dm/4YbG3Rabm2c7+jturoRVofTF9UnWKdz5r7gTnRUQhjt6ywhfcfPrF9zMBEhvHiydAPzAveo3Yf3+xE1MOMFJuBPotwzeS652TYGO/PFZk8AZnCuVTxOMEf2wc7t/G5kzz33LjnyHA+Z72J4beQp8t9eR9eHxo06xykXHI4W0uoAYOHH3KU7PQg+GoBpLyJA9Bd4R33G/ZAG/cPMbVuw5DSzc+ZSTzwz92zLxUXDjsy/yejjrqP9furyHgO18onldz80hn8lBjvINt+kOgFmPMQdLfeKq111wVRvsG5BehLU1Pu+4n3xyXtVLerw+8Yr7JVgxS6IBS1Zz+drAnccpsrQQefc+ErYjW/80DXJQP2w7kF9Rl3Z0nAzA0p10wnLZixuUPZ/02PYsFfhHbWBMO/JZRYJW+DnfbbSOTTf+Ic0UADMCo0mfinjONKVpy9mJBouRjyLaC24+IlY57mkQ7mh6JaMZfT01hYK+bziM4U3QEYeXjDb9sh2f3+C49z2YRutOxIcVQE/RytF7n16sNNn1AxjMLGJ6XcFf68sDnzvwF8f4cJYLtw9RXQR0Ank7hxp3nawW3sdDp9+ctPezcJd+a7rcMwZ3dHxWWfPC6IFMReiszAK9Y3ScrOOV0sBJ2VmpfWHaOZb8KehHhCMzyQCLbIyQ+SaYx+8vU5dYtHNaSE5pTznZK/p8POoMfBTGVp8ReLzl5YE7+5rI72cYzBr3i9IqEu6IR2U6/STOKwEwClhTsVQUfWQ+y6g9+3vw2tp1p+/DtsLvi/u8yB24m0XYaX12NGyAT9zqx+QtjLYoLcsRv9VtVkH64RgfQzXM77e8kvpMmYbh9tdW/PiMYcnC/laP8gwlZpB1RzsclzKHq4bjL7hll4gv7gSuXjzlS1GfKRF6t2fOcRM3AI1NaXtosRWXf99PBzI3OmHUCaKc189q+huDddv0un1SNSPdnnJL3ffc0h7di2oCG3eaLi3cW+jCzft7wYzoKqe2cWtOhcZNh+5ZmTIJc4yl1AffTqvRMwXWRxv9C7808zTX6KTh9pWI5xLrEWznHvSxPjPW/eyFggDmNOTCXUbxqLONIY+ZUu6Nf+n7337i7r6X3tYz+gNpdnKpjWlTKcfWu4U7mDbupedjqFcL0F7twwJ4+LNYdJwuv7hivQDGmYeOjl4ErPQkRmGEDOBzdb+yBveUqf+2M9sR5SoG11vX94pAoBeTWeQbQmRk9XbVflgW1ULv4OgvbSET66g5TR23MT5weB1gp5Oiwe/n92cYRePtZeWtGFqa7BHfxp6nqfdpWkaeo0edKfrydedJaOVonN+z3IXjlr60vGPIdA1NLYLtjVQTd/Z31zVHl3zOg1rm1AW4A7/IvXOLAkYPa7W+J2srf3zaSGmr/wG369IYBozga79XRsCsKlTX6IyhHWQ7DJ6NeWBn88adKsJGAsaHxzAZwt19PrOYs+pqL/f2VwIook/j6B78zyZknCfhC7OiHVM8GGxGXMx+P3qvGbM/836P4E+BPpa5W7u9LDY6uil1gzE3oL0JIO05nn0oEe+Pz3C+3v/bgiI5aw0N2tDmXgvDbZmcalL3X+/eXbNBE/cefgUYIaO3FYGH/XT24DUgw+51g2UMrNk8T5UyR/DgB3FvIyz9qgjfGaENu4T79Juu5170M36ewNXOvXGvOtSg5Q13T5fTQc1CbTQkf0v8YEvruS9JD2anxZuHjuvv1Z5wr+/oPOPMhkQrnysXH57CKYQTvKe6lmr2dI9xUWPYVuI+FUrQ370fmZT++4tSKgx41Lbr/P0xlbSe/zfcnikt3I8hxiD/0z3se+RYgFmPycbNMeljOGTPDtyNwd/n0f29OePAnGqDsTemXDUcNb7kbgt6ZuNuR8HPyijc8XgtZMhq4R4f31W6HI+KkMYTrGlEp9WznayhldjrQaF18Rfu82cPx5zexlo0/8RdMyyefepe08Xu0Nozx872fultXMCd9cJLAIk1Zk2LOI/IaEbkv+s2Kue7wRx9Ilg1er4Yb7J2JbCoPhyPRxlbpPWWpj6cgaeqWPf/B9zKvOq6cLewHg4sUVFo8yWrbhOtoMPQYz6yi3HhfQK+z+OpwDkVwvsbWRkdDn8azx/R/xfu7mcGBMzrno084oMZ4Rtfd83B6Rsp98ZtBvgoJIa1Ybj3UEI/lp7Y93PHcn+XDyf19vgLbjfoNPp0r/FSbTlPYHtztnMl7vVsOcWrN9O2t3k9l1LMuZvJFVncucsbinn+k8DfDNi7fPHAI+oaCGPSY9OW1yPG/dAzv3E/8Y/j7nx8rN+3g1he/WGQv/pimzQw+/eCe47V+dVLtNo0sZ9tSM4n8R7z56gHvUVTzGceuD26ecBZtOTGvDDJUePpyGiQ+xON63k2qz87Z3TYb//pcraZHNEchtvupbwKdz74WfikA4uuEST43AvPt/4BNtx6GG31aTwzeWeeeZDDbU4vjc+7t3x4V96n21ld9SGGAX9Nd0xxRnGUQXaPnaOd1XA+RnvYfeac0h3Wa+q6o9dRrFGMc2f3KFxR0V4MUdfNif3AfT4r6r3iXvh/RKuN29zgkqnhdmP0th/OiNH7bgN84Ebf98ZHeF/dPqeB82E8W/9ecNMx8HutKaFjez6j9P2Vp2/7eCzYbPre9HwF0BBt69baFPZs18CJTm8X5mhiYHlfw8NH8kmHOfnvA0TYVnQBcpD23SN4XfN2lDDGjIpFLPfEDmAUwELAu3hoe/C30lqFuwmxyBsubhoaK+UbN2lYFWTdQjrN0Y6IYveNFHnRzBkWzXfHv+PebbwO13qKlMporrfIsinLckJH+pae24zJQylfploVdHw8PMbOlIU5qIhZaC2sPP+E+5d+417XXoPRm+GvdUWFIVSwfqv9vOic4x5Z38btcmKTdo9Y2/rSWwjc8T5xn1lAYEyBb8frbT+K0O44n/Zd65PNy+8UpxFZA/GMjqjo9DYuHWnkAouETgvXCsd8NEHjed3/UBEnR+SynyNqn+t9lBr727ijf7KftyLTawrr3tJ5C1PiihRZjoKp38iAXnD7WLUwdxQEnoybCtARith95uPcmxvDzyxwy5o8sShYyuuOb8jD5e38LppfcQON4w33znyCp2O9ZXp0pi+BsXjsBpbS15f+Bm/jP+C+Tc/fnZjj7jVAXo+bn57SnQ7kiZuObMtu6bRwkxU3vriReZU3UkQ4gPYYPuzh8I6D3rgZOwQfMKexGKOpLzfWHYXp5VP3dlaRxtuKSBW5tIjIva1HtFy/AzgLgjhuq744LaW2whR8DY8Gw0wxAMA3jOlWw70jxsiSis9DoVPyOl4AACAASURBVEuJS07NjrWQS9HkxYGacty3yQcQzlJ/0fDEbYBcZpkN88fQSDzyrGVP2Qo36eUir43bJTDC4g/cACJxm17OQUYi7q3jjoMyoNOirtI2zpqZNkbXa9JjRBI37QU1xZp04dTDoq143OtBPcAZnRt3tZ9Gw8O203EHcF349l05Gwdm+uOe35U4D8OaZC6qsZV6I3oA7+sugJHWDod7hJRJOBgC70NUpnFog1MCemeGYL55WNhzRhMXxqSvAzDFpvCE2/kYJr9yMg/c7kDaCcf16Uiv5biQ8FVD8dQ7evVriAYqNSnPl+0zUzHB4SPuOjnJ5CijMCym4CO1tgj1+OwsgGiJW/Wcq+VHfK+4IfqPPpIe/viBW4Rm4867r+ddXdA5c2i3HKY5gg5Oqyb2quO1iC2euHtCoBbGld74Ce1SG5T9ZfVTLzhyvjidkdkLMgt33HZc4ih2cov6ju7q3LygRTT5IPNSIcJ/eDetJIOM7ujxikwKEU2PnMQj0vIeOg1XSvc2vivzMCmBZorjBiwaVDvDoeTAAcc92vOf/egTN1b/jtskNaDttQj+rCm9jIq4Se61vrP+4xduv2wrBCticbm/Mkk5Rms3jV53/APE2qNTMh4ZEhcquRNeuMMdZNHzqFU9xv40EjrYpkHRlsZXOMdrU4b+7VWhwAiSD9VwfjfuzuKo/zGeE72O2756FHCXgz33rdqhRg1OX+I716UTsys6I0UbAD10zxX38mEWh+47Mc72c0Ykyu/vI992hJ0RZ6Ge4J0Z9sTDf+Q6h0C4fROTt2djT5JfGZPG+MR93+aESH8NoZSBLIV9/L1wj+zE7hm4F30yrjaqXiFJmXDWYkqg/Vzjbnn/Abikkorcwu0FVle8zVPvcON+w7dksRwLg9fxVQE3qj6MtvhB/iySfPjNGRPVTKr4Go4LQCrb84J6Z9MqFO/gApiOwPj1H3C/yTtwsgl8njJz+yWHA6MPFkbHNdnWjbPk/VzVrtPjPa3gpXcpJtyhIK52SDIupmmdekU8laQrz2VsqMWjtx8cs7y9G+uvRSR5A9dHCqCXsmgoRDpOKBjnEASq/mIe3A3WFchwkLbTpy9gcqU/HRyncq12gbyZKqPvf5tBGM4QrTiSRxkGAKWoy0ifWVcA+MOcYfBoA/FcKmpDT27mm7hXuPR7Bm47RZu4LxZ6lxMcvCGtKb7GwE09EQD0e3YTnK0LHadodI8ZBGYQde2KRVsaPxY+6dniQTnbPrSosgsOA7yu8C+4faaDGZgwRvcdVlM6786tzAQfo222xzZ6SfsJLAwqVQzw6jKNtJnWF4jaKr95g3vzBdo/ZqyagbA2e1rMpue8T6bMb44C3d7R7QIWtr8E53dmS/3uEKNX015d0O3syrxs3uidpF0A/rf3qR7ce+aAfHLjXFNvwwHZc7FwR8/uHAdZBhD1u8bQlGvq+X7DVdP2WEuSN3Q0XtHdO3Vve96cu+heuoAbuG3KW/+u9Rym0/K/jbbMWz33WH5uOnzD3UX1PYOWTXJm4y7ZM5N+nilaAdCc1PjU89pRLIdCpx5Gk3/McVjGLNzRe0yOLnz0nNez2qn8KEovvZ3y7tmtS/hGimVGcpuiu/ex5bleJU5/VlmBzaykgzl9alfpZUUcGfl2EoMQw7gM1VI6n1pNfV9/RaBf9ty0j5kgU2yP2nRIOz2lsbZhNb0bN+I6i46AhZsKtTOC+bvjVvQoHvsipnbUC7/za+Mu7JLvQ+lWWxqf32fZvpSduN0RXAPvxt3ZW2Fl8BrGc2jymZHGkM0Dydnxsj3/547PjI/DteEAV1uJYyuSt+Nug8Z1yTHQsfkZoO/6Tp7FwH26d/kz6FMXiNtlZYHqbamD49bfF3BnfhGRvRHFT8qix6vf3fuzC93mpaOdhvF6PSVZV3SryrcvQ02+Zs6jAVvx9JwM2OM/cElu9ixCSn0QiPm+h/HeBAcGOTumrJmCLLR9YUecwa0it6b7rOLPOfnWZY57zdE8ajP3C246a/QZIfxUeplhCsQj8D27GfKfGEatB0Dss0MtG9DsRV0YuEuufQq3Z2gVXHyrdhnK+dWvucMgm2gMZInro/1shRBuvlag9ZQaM/dNjV2dmEHlP+KmA4/nYrDW/Y2bW/7bkTW/2ITPXNB2mUUDfvCOmGPZtp+7oSZ9ycEV8c2/v/IV+SReTHAlMuJiOwX7QwfaMMV6M6B9XDvaOEfKlBgHqooh08SnklNhLC2nkgLIe22ce3zCmvPC58s26mXEx3d4ZCl6rPbyrPg7GneK/ns+2fjA7TTNZxM5X1CTzj2LWgE8XvWQL/xyujN/4zY6/fhAXBf6VQakwYJBOs8s+v+rYyb9Sw+Im0O2UR+gU5jaxOcVClfdjIuk/n/jpj151uEO0HF7BvOW2QzcDDDodkCHYzUXr4UlTBcn9uUg8zqp/0vHxqxBANB/b0PnvU6UAPtY0pRyALcIt70ggLGsmusfdrQdGJx5cYpo5XFnqpXzGfbN7ER/3830jRvtHLfC9LiZVXVv1/FZ347LjSk6jf133GzH7tfv1m96//+Ce9BruHPhNiN1PoQK47PvVgELLhu3hi2fScIDt7Wvek3Y71sepIM4vXGrU8hhuXM03IsrGzc27oEz19/LmKOHa++4d+dX4728uIvJW7XjTqyujbKBno1rFoDMU2+lYvU4MMFo7OQrPlM/km1nTdU58OF83VGg73mNHmy8x+fdxsSh/pFdf3kUH312xPs9PyWssPUUxH3/oVd8Eit/nn61QQfbk1d/sft1g3da2MW9Ly1eWTQaxehuTyn/o53lmOqeWDTlvVf4psnb6ySMbGl/G9yrhoCPLC/FL/7dhvvkydAR8v52hd88JRE7UPA66byGbDP/8KyPBTScZAZnuPGGO0zOOzgPOI57GEz/pL7B5K1rTicfWbM4u64i3Edvj23/xTUKIWFEjMpvGjHmpWR0jBzuTI4guvJdw4h7ra13hhsjtdY9vOCy6hXDa7PPa/D+cZ4mDaoMyWcMGvfcrj5SyEk44vpY9CB29+Rx2ryXF28K678zIxnF3TUse0yN/prCU8rpDtRwLyxyLs4LsS26GZzpuMm7kvceUjxmipxuwyP28UVG9bzJJpS+80LX2lpvXZcNGw3pMetA3G5YPuS29CeeBUnx1zPK+8Yz+puOFi9jYHPcuXCzD/LtsvYWnK3vsu/FI/s3hlmYbZ0h24XAld/xpTx2dzDXPqDGfrGeGb9gGsUN7oIfh7C6ku/xGdIctl83Rg5ch8lNVu2clIK/MBV23ce3wr09uT0jHIY7MO7vRTGMNIV7G7ZqL7zHi35phrpqRo8xMiPZ3U70jf7XjymUakbG45F+P/GNlrJPSGtMPIq/20kFnpKVajk+++bYjBZmeOO7XLiXnjpW6XTacyEnmuNwmDnsFL6VoZzrn0F/DCfP59mvT6m/4A6g60at/36841E/6utse/AL+zodz1UqWHTyZd9WO4nq42wkG2kYrGHogfG9g/coOopRw9VBG7G8TmDTPBvfo215YzNSKcVca6AG3QHJ2V04C2P4chXHDcO6cG/ntJXoBffJFD7IYSjZNJH+R9FwDv/O6xWMLis2q8L9oLUcUPaiMeHGohnR95kzODy2dQAuEypRKajXogIfyeMdd1ibRu/GXW0MPtm05G/cLm86vqv7luM1eUcaz3JuTVCmStzk1DzsJuKDMT3szn/QEs1PZcMv/IDdooCBdqz68vTPrfyP/ULizzVx6z4JculiDHkjz0uGzsnJ8OPh0R0NQ9iK5m2bQPR8K20bpz8TAtrZ3tty7OxpOhNqlBGAi4vSV6uZNzXv6ivW5lkG5L05xT09qV+9GOeROGsl4qHpvE0+R/8bdxAfbPl7KdbhS0xe3v8s3GzSV+kd+n2VpO8q7g1q5Ikr1Zu8+avRj47EJziGXhPR2wAskIDRkkuR62wO2DZx4XbnXLzKv3ZopkiNezkOo9Wd13gFwnBcanDqqnCH6cfcyOXOeXxecQf4tnX1GgG9cc1f9ZnZpKyMurG0o5kx2nVjzTr+ytjyt7zjc5Xrz/KoVIKV2saOMOrYU+N7dubM2sQQTP19xkR1TwC+cOkI5jPu5zPw6DXm6pcje/xN8lz5nfAYfbTAq63BiznPruKSGd2Ymhq4P9X0JeflfAp/KbQC84WhrGUovhCpebfge/R8y2r49Ijihnsw757sGsEjJwle0yEuyi4bt/bcXMWHwQtz4urmBffIjHmbF1xJj+nlAY2xXFzNiHn1880h+MeKx9fkr+OOwMAYCJu9wDtuc3TP81vedP78G7iNztE+tr7MYW9m1grOnTIpvT9Ko/QmOSee0KGwEpRNVXnKaallGhMG8Rof8vZY9ySQf81cthNDAwcTRpYgRXLGGG0U7i/cXKI8IiudyGW0pzmKe9LwhhvtMKasjXfboXkKT8fuig9XgO38Xwy+orgfK9DL7/ecvaiuNg335ov6MEdJpxuTB9ZqO4i3wLNrEK+4qUsu7wH64eDDgg1veeJme+ZohhG6U6HsBAoKgswO9jqWiC7++4yg417D+xav67fJfuuUYfRXdQwz1b2O5TjSa9wwtJZrxMudaHzLFGkT/67YczwLY4Q5FI/YAn6YNneCvqVS6Os+DnOB+78xRPkX3NUWMy7tXtwR1CMboxQAH6+PYq7jZvs7ysens5qAOQj/EMPTMOfKV6vMZz6f5XSf1hRcUKb56NOczmOY57j5O3E7PRZMBu5AXN92FqJzG8qOoC+4NX14r0da+X04ohW0jyyC/VI/2PYTtweFNl6fCfJNjR5Io5b7L33m92+4Zy3hIe/XvUhF4zh1a+uPG87o9/DoygJ4GPC2VuI20C2EBFrRVZOgh+91Cc9xnBWpXqOVR21zTvqO7UylmXs5iv6RMfAZe07KtKa6Emu5dLZSFe4H7Qd4Y7v/1vNWGR/RCnhLD9+HhS+f1yk6x/uS2bjc3EASNrXdRte4/6az3RkMlhxKp5RCiwZmlHNNTXpmNqLlD/p/4B7vy8jND6t/uF7cd99bvNEKTTmI6kfDquVIBu6E3lI+ssGFO2jsjhurrf79eQK9YfB+Bhbyxes+LePzdd/7wF3Pf8ecMTMBT0GHAUP3itkeCSoSphvaKJjxefOo9V2455Vy1VSWmJDqQwwRPe5IyDMfK8d8bkR7HMHy4YciOBaAJzY1bptq3NmVf3wsWxEoLbr7lN7B7YCs3R/8nJkZDAehELcTZRnPwN1FW2YLPIFJxbh7G+ULfcQ3Mo7Tb+5nNm4O5XxoMgxq4aZ8fBbmIf+Xw55GIFq4swvAnV0uh/hreJT3mFnRlLIHi2yaJu6lr4XvuV7U6Y/+c9OVjpu8wwxgbks+Kii812uVtK5NprbHEsGshNsMwwuSBjNS8Saio9xewIOTGq4hAXjOsBTT6gbDGCpSrbMkHkuXl7AfyqRmo53QwL0cxWBG4d7ORUMQX6TWSpRSdIui7iCSfdi/R8pKg/mBe2F8yHs4H7afUnrPGHLT50VEfVJ05M5qmKr7vfvxkYk4XV7v4ve9AOu5qM4wSjeBifuy7wnrg/R7crYKBoIHZPa/hgjepz4+vfoig36wf45i9A1oI+bOtn85SJh+bl06/M078xx+M+htDzaZ3MztgLemFl05NQTY9wCPV/NlgicTBA/SUZ9XGZT51D13PlKzPtvhfQkxjWJ/qPx4V64xVfUWTQAdoItE+PtidY/NMsTBkcKNppsNvkTriEDeafJqPo7XIzzG/hv3Upw33DR6T2llWPP50CwQaXeZrL+zF2xxEVQXkE13XJ9GEfEXbhi9Td+YORpBxR14d//KP0F/0nFEE33fwN08TTpVcAqV7tEzzNaN57Bk4vIVrr0uxXF/mu9m/ON83K2fO4tjxndd8SWmpudu4t3P5/P4LXjhz5kruqzhRBkRv59evJ0D5WUH9K6xbR8yaoosxapTuiTApn9439exoU8XlRCzXoa7mK5TvgfuqIA4vbbaCBNmonBbZB/Mc4fUhtCLhlYRK7jqtHgnHprQ31LmN9xD4Vl7CZP3ypREgyuy78acSnyO5ks9/xwWeLrcPB5bqX/h5vBO+mH1tJ15Lacysdtz1N1cGAPjbeavuEEoRyfGWbBY9Izh02U4Nq1RbLkWXjQfRqDG6GcObz1IuU2GnDrtqJd7dziXAzDzmoxkI+DGKh+GNNj2ksA5zo6GVt5KxnYv4jh+cwpMMbeSqh9SDXSaVZEneow8cJkBbdw8Uv+tb+EeypLdr2U8jGyd8azoYbgbqykGMb4aZ93GsbVkwKnfF9wm63fcvl8AIyg0bsvuAMBOaSIfxBXHnQBT7aMW24HtaNc87xOfAC3cStOjIvh5kpUIOdad/l3+wJ3j56yD1EuhiFsBYOJueZlzj1iOxzH73433kNoBerDHZ5vqtQRptDRu159b9zXn/wV36eXXj+XiMzrcox7SlJKP32Y60oZjl2jA/kWv2dAFMVseeSkzvH9Pnwaw6F/Ne3e/HT01pecvYTZPz/eONFg3nI2RQpiKeSickVbBZg0vTjPXC+7ByPPT8fs+Haa4iWHEE/c1jO+Jezujbmec+GQR90lnobeI2I5i4h7Xf+EeNJ1ruQqrukVOjN9FX/c25VBhuF/k/fYZ608ctwWMRzBL9blXqyLWsyBtptukNxPteF4mBPy+13bJi5KpLj/t+wE7LnzR3KuLvexY4+kiwl3FXqM+/UL0KUxrJdhjJV5A6WXTaoy6ohv2oYTRMhWVCuHXPYU1JhpDx5DlF+6gt3fmLsOhA8iJ253SpPPNTtKq6K5A/vxSev4+XoyxlDLtmrUnisbw7ZzRyejjY1ztSZHQ0f1s2ox5vc/Fro/Mgrz0AOOGU3/S2Q9jK7l4lutDVd33posexEpX1OfGjdFG3+Ns9+9j/Ayekr/qCz/12ttSBuU2ZLqoYTltauLmVghlumu43hsfJ25+1rtOOzJ3KkOlvWeknNwqb1/EW0X2EXV3JPZxKBXJX3yiR5fnVvSgwlSfeib7fsCUNADfT7JwG6ELNzH52g3SQuZWEzLQfpPZwC0BWlsUtk3dubOzxptX5hAf+1wS6JdaWH/6ux1yy5VOuWRahxN3AKr1FjDa3EEANuTbuzPZz+z7yQvHueThfLAh3uNcDQB6U5ju3224zBfutDqNnic/MHFzCHvfcoajoCoH1k6h73kLfps39ruCL9pZSh/QPMSenCgnQH1O6jHttXAPzGjbqjUnc+p0EOvMZVRfjdnv8kbuzQmqjKXt3qOkG139vRdE6ZVwUFvYbckgMe4dG34AdCq3YLuQ9PcLbvJFkbQVd9J1kYIXWtGCdkUY2ch0dq9FP6d+y/ExhfemmMsBY2HfTFK1/DZ6YYoMcGdxOLYH7k2307YdxMo6xvW3hX3OJ5j89ocGtHEP6qxdyqhwM8MpvsbFfl3e1o7REUDzUHpFHQ/DwQc8k6jvc+uHZxwvEB64/cvpVN6K+UC9N6R3pVmEMaARV2WGq2cbM83MazGthiTxy8gRI0sewAJgqtuLYwYRaOMxwZei9ilWe+WbbYN+NeiVjvr3Plbcyj0wGn2jfbtPQ5kZfaaNhJCO6LgjmOEeq1N3WjyKXU6H4R7KWJFf2dmidTxv9LtOLdwU65gyXZ/ego9hmOKZK7zjHs3FS9ulb8nzQKzdjdsKk8+hj+Omjm6+AG+4EWFBMfo9PQHwnaZqX454HVfw5mSHPlMO6HvK0H7jnn0i6qgFBL48oYcRIZWq9kfTM8Zs/3HapGFR/D6vvoTlgq9eUyCus1SaQ4vsabrngcJ0ND5vfHqPy6rzMZ/wVFG4H8tod7R2pegoR9x7pqdxb6Gg//ZIMvox3MhFR/MtRLfjrvdGVb3BRZWZvWr2+lTAu5dCoce6I9OhA5tGMo42+GH0b87jMSTx5+kLRpq92l5GEcqk6gRz4+bArbT6heY33FtXq0j8XIdkfPLh1S/cu2aR/bzvyerm3xy4H35EeWfTFpy9QuPGbmM7nG3bPDcF+b3//sF1/Reen2XMjzR2Cjnp/bGMTFVaUuDF06PUYJqWifTdq+zHq9/F6DPVyDcmPWk6DsfaXtE573/6+9i4lrfeuIfOVgZzOl2PLGcg8qIji9U3+nN1W+FKdJQ4ypEmbIl6MSFhe1I4JDxcatxU1gddhvFRM1r8yJcMhLLmc2HZ2+jvqRPdxcaNWffBDcAN/xjIYY2377jxjlv9G7YVxCZ2Osh5spXWIFHWgYl71W5m3+x31n6OXtvxh2ORY2c4PTOU4hs14dhJtfmQsWF86dt/HtIDV1wRfTMf3GO5aiqmYJMe2ot9PjarMW74WGtEaGdWC3hGsUDXPep7nnvpuGO1bW3F9em/RwpdCpD/jrvvbeUYy3Yd9xV8dRN8O/NcC0C81e6uu6B4MfgGXNfXIknMZyPW/XYuBNt7iyqS3VrkdVpYuGG4f9UL+JzJw0n+4ZzHLNnAAmg3qlpP6FT6iOJz8+vI23A/MkTX1xfc4bypu4dzmPUF3zj5GIKTcQ+dWnbwYisnS5z3xxvu+ik9HwVR79dqbANDta8AVzSbvCMQ34jYnMIQnlLDp7HrmLYiUEMVq4hvxdgvO9ECLDKagn3wltOz/dM9Jn3+uRTGsH4BsBzDiFJudI7beXi+G6ndA3d5dvf+ZLrgEzcj7jUgn2Zn5Jv1isaotDXJQ67ka0y5Tl3qdt1Bm5EO2my/B7MEys1x29h2Onz2lE18entl9uU0FQHBvs5PuTUZPXUM4JmXM3vxTHPTNHm7DZv6u3f8xlLGXl2Mx7Pzi+5vZGHi1RQHot5w51nVcnZJeYOnjVUDyVm7MB7bgi3x1wPxdNRj9GA1lqIxrz7gdUcDNlLrDfJveNcR2SWk1BZnCT8BT1XHsfn7I0dx970WBXqrNC/zu3KEdBSUwJboI60kbotisRxG8qwHIjJPbLjHlnQqw8a9P3IUdd9N3L1NnFnM8SPZimBGSKMeaEfau6LLcBAdHbloqw8L7j6eezeKnh2Zc9WWVnTTGFp6wX74TtVugys/53Jk/5FP3AMzDdKcHBlv8j6BqnDbFHjQaS0epkdmNzTT3+csI5oW4r6p1396TjJ/4G7nQk2cXUzPM5eb75kaZjAMVvO1Dm0Dg4/xjbhiRIg888lnQc7yNuKWvXTGI7WKZYzaBWJPLdpY2ESAGeWXh80b1+VjxdD1HtdZO35NaaVHkX12Iw3ap33dMZyInfgrHvVKvOfYUkRjKKlF6WexynFf1sSN67JTozlH7mJZuE9rNuwaQ8PPVGSTZS+nnnyvPKXaqcwl6tzIXzMy7LvTiPpqR7rGMA4UzrsWEbljIj/dalz/Ejvr0TL2zXMNMaLk+cQt3VlynPLugHW4xFoami7x1vne8GfgtZrEwI35bAW7Q14+5Mz+N245YGL04KegvHGfe75ADCU5RnBZd41M6Zc2MtErVwZRx/73CKa84dtU21as0aN9V8zW5pjVxhzDO0NtlmAYy8vhpcK/xnslBPUdl5aIjz0SVJbHEGZPrRZuH3dkzlWqAzcWPmt/92Vt5zDChKf86c/7sCrtKD3DPc+78Owz1fbAVdnJG2lPXhBXok/YLsfyNvYfNGwD8sVyx4AUm4CWuQ2Dmj/X2TXLuyOgzXKamXPcmLjlSHzIkkYPf7fnvC4yhiUxWinif+DOV0fRKzIxdR1um7UR0vqdPGefdJDprwLwhv2BnlHIsXoxGkgpwtv7FBqgRdAk4Tb95ESL2c4xy1Cwb3l5Vu1NpdKmKsl09UMh2mrUtNPDj3O82plgRQZP1wduDOOcU6zrnvHxqvpSuscsSvcxcJPl/csLbvKRdBA3eeiGW7j9gFnLHvwefRtAH3izDMpvNzmOlb1jaHgvjIc/cc19Ix04l3MeYX0QiMfq48Ff4r6sicWX4UDRgcanqI2m2cwLbtjU/A/cRy9ue971z2mk3QbObmKTmeMez4jW7KrLazQwxpbxjLHM27hYTE+7j3UK3gNwmNIrLK8aK/HaJUH1GMqibVgEkiLZcOcRmaLbiXjHO8GLroPbv7LZo1eBvOMOOlfPiDZuOiOwjtDN9/f97Gnbo+JyHuSX+Ob4jC7j00/ceMPt3xlu3YeyUfY1ZfiOe8mbqyPlyJczHDxpgrn2omcrHqwR7XtDZcig/d/E9IrbHAGHCOG4L2I2+RZW6sHETfpfcJMnOQjS/b2WyLHSbpczkSzecJ8OvpBgdnSGhNeNcmoMTaSGIdk/B1NjUBtV8T0017bnETUAhBlTQt76kFmMlPA3fRR6r7/vBORu+sXFbez8vb5L8mEZue7Bei7R7/po7D2GTqXISgOVLfieASiSNJmVoLojzOxNZ+WMtFHI2mk7ezeaMFonHrIqir9muKMG4PLo3/sdJ47nPNsy/DfcNCQCtKg/Iny1EV0UlbNLvuCqonA6D7pN6TUzFXcwjynJwt03LNzc1p96bui0fBPp+jfcO8O7ukvKDiVvD0Z5azFa64035cPkHkE4bs20XZ/8orcNog0vOyK+OgLrcaXQXUDx8xmmUQbSlvoaapEREni/NOjul+jKi7/VQnyBic1CGIZNW085Erod9MP0j9S6ohjzX3EPZ9TX6O76ntJFEHc5F7zhzolbcskWZfYJXL0ZiEVZ4l7TalHO2x0YI2S1ee75s3tg7QIAFd9xVwu61rj9sJoWkZ3HcBmNL7jPndRVyqkmFQ0LpxnPjcehDPo8vX+oeOHRbBeH2l7knsb7ituH6GLBxu0ZIgy32SCAiKpV5KEnld28yJsZ3bUL+tuefdUq9B1Pus+843vUs+fmVeEvFAGU0ALc/tz9cQqmOz0iPLMpOreifh4F5vDjxVEMp9Ke/vy06v7IghywR3Uoc4Ew+IL0ZpCfMUDFUhpsii+hmoLvT7D99p8gjz3FfGK3GKXowfZhPAAAIABJREFUtHHfgGYMeHf2j6CDtENcOJMSYbgph3IewkSlnelwr+FIXCMzoayN/uKbCow02kcUJtaQcr4OlzQ8mGt65MgeDjtKLzdu6gmzy6ARyHHB5IYMOf7jpzygcTexWqrn+nrPmEwHOT4B4Hbc6/6NG2+4c+DGeGWmOcUK/uTtY+ZL7yMmRJ9NPL9+zwOf5fWoqLUSLu2FO5iLcWZkOAwK7WtAe6lwI3WqPIpFe1HPagbRL+sVBnNT/RUr645WxK6l+qwOjHmNe3h0NJPbOAEuQuvoxyj1MluzCmCgQlY7xrSFkVN5K2KTGEUTmHxqOZnkQ3pocIb76msxeBwTt9PHIY8Kv6HoPmsAT4cG8n/gbp48f+9MhsHHMwFSfqIphgMYhrvYqnpJFo/7CzBTbsyk3YKJ/t0t78Tky5B5ZTfE7Y7U79Pv00Gk4452kD4HphqNywd0kPXbGMre+pWLKaczObL9xnVlK8oSULKhE9VchTvy2Jy2Uq5uIxAV7ANueC2C6fWbjJQRtgFYRbm87fnzFgPSTo86TvRiXiDwioARmJvcTCETgA5racfWDo96wP7uTqErQ3vi1k4FjINfH2szDDfxpX3PYZor0X2bQ85ak9Jz6sEIK9xb3jaceLyMmbrUfE05rsYG74/3e1YZ1BWqyN1ct7H2K27jicbVldkM3FrNaj6M06ByCg796FlSf6pVDUVNx+mMHeGRZV0tPknu1U7HQBr03WRkZ9qpwNlDCW0Mw43MHsJyyHKVzgm35F24r+0kjQHlrDqsvOOmLnzl0YrIjrrVYKVBQQ99+eal+t48tyLaNT1amoCbFO+Mu+3qCXo49dZOwB3GcPwJpU+HDl8+a06Bfdq4W46d3+ndHsA52MQXDAHMSui5E5Dz8m56GCJkLS7xzMeLl5TX3IHrpiktjrALN6PO2ejECIN2TN6G4abu9/ibxnZ31jl4mJLPjFLNz1T0rbaTU4gwXXHcNMaNm44I0i0ga7n/EzdM3t7/oSvUbx/QU/dage/oTDsdLyjSDn7jNk2L6POHstv0Q2qoJMKrny3zsaiKMq1gcL7pWSSgDV8KiIlbcq8sUzWQwu08ED/jqnUWtiWWoorso+7mW6buySwZOMdOvT6hn7FpnLp0w1bBlaPwLOMUN0+mMFJaATXj9aPK+JJhOYAucj4q/tlvMJdHr4LRGc284SZDbWkyGbrDVjLCk/SzApQvQj63WF2l+Hi8vV1nes+UuZR6Or061Vx/J3rcXfgq5GT+0/yoKBW8F+gjAhI4K1ZJhp+AVfKKotmwBxK9JbyC95B3diDxUAgaUuGy9EBHIGiox3gY8PUnffiw99cylGckzQo2t+1EBvj2NWYcHSdu65PYz88AENdHWTZfttVD0TM70g7FHLh46LjppJ5OeM4gZuMeAf0Ft60MPTj+tDYlGLDT9Fk681fH6tXZBvR4ngEcp/AxomMar47TQysrGURZ6DxOshRLkD72nU4lroDSblcUjvdGKCczumbSU36uJB2V5PYBhLKo/yluRiV+P4O1p/Pc1DVmSu4XhW6uz8jk43vhtsjpC7SYJaB/6roiJZ2j4c56grsdqaQdKs2Bzdmdw8bi7eWzS1PePWTyttLaDGNgZ5P5Jm+siByWXcwby9kc3Wh52TRsBEJHNTjuNvRJcwwySbeWp9c9RkAdsHwtynhf60/jtiXndY1Tse6az/+ZEX5W08S98ts0/dWsE/WOuNuZRdThNx2gmhmJxMWDVJJiaUOiYWa0sRD4WVdvxuHjYyorvZ0qy1Fbu92xdKRLE67Hbw5xHNRImVVI5bWlRPZ6I7Yd13fQcO6j1y+WxGT+IVthCj692JkHnZk5nbZgffeOu+shwpFdHG3cEqbxm9fN6TFqDtyXmNvytmlB4Z48HENMOewX3HLgHBZ5gdPw3aXcRY/Ll4ToMGHHTNzj3v70WpeY31/ND2zcxMjIyz6z9fMVd13rKVwMZ966QJbfp95WuDU1+oY70tp0m3Ed+I1b0/vRTp3It2ydt1/kX2Se8yFOP/VI4jgD3urE0RmEq5qlYx5icRtzWDD5MyW+Z7+ATjqi7+6TitlFWk3kDFeacdWnCV6ANQcNE2R5ekYXxz0C2cZN60lheeKWKoG1j063XRFYxDL+bdzMRMygj5J7dvIvuOWguChsvdgpMRxMU45+fuBufh9ys3WDXSEmbmFh210Ipm4UMDlp0eI1BgWi5h8kQ+J44bOGw0Z/ppHVmQxAPgU8lPipeeMEPVvfwJWYY93KMPqiLfoKFI6Mp3JCs9NuirhNr0fhuvnjSxyk7+ltmS0rg29eAMCX3rEjdOhh53NfO+m5vFMJJpcCeQQ8rMkyULLEvfue+qlx34Gp/w74WW/GUlHW76CS83dXDvv5P8WdgM4hBSZuCcwfCt03dk0qOnl078ei1kTEC090XiMd3d3z/E3nxCDcVFAaJf92m9oMFpIAKI+r5vB1dN1SZDkUyNg5O3WcwgvuiFMfixX5xunwTfdrZmBH0o1MMg3Y+N14FPGEXmdzHjWZ2XHPWLRRChtJsYKl6mSK7nzICuMkx7Kvjr2lZ1w7MbKJpuD8XkaetR6HtStlcIHNuoGk9NwMUXaWiPOSIa0ekyObWtTCD/BofC1nrfs5jNBUY8yIozcwDSHSi2UrEMfPrBPQkMXEXAtGrh7Xq70pzAM8u99huLWLVI7MFEAehVNVPQsg3NGGXdy27lNR0QiuGHKPa3zIo+VRNJvJyOb79WnHko6b6asUJ1c/VJG/pit+4Iax6zrPHCo7m0nKxNOwNNzxL7jt+zZYRsGja0dhWy+veMNdooc5EhWnWcMynXvox3Rw9HvNj6a5Z3Lsb0In7o+tW5Id3eqh61b9HMDaQRzaL+KO0nkeLUCwaxmBjJdBhUVqk62/t0X6FdAEh2JpOe10msHTvW0hEQLzRSjVESMaAUj4Hs2i06eWg77nctMxztTjxwh6BqJyChYsQaYASB9CtDB7L0hFJhVuFiO9LfSKyFhZQphjOY6Bx9yPfKCh+uyOhAH0LMoK49XH80AgM4KxfB247z/jH1r5qh8tMuIzKi6XOxX/v9aCrfnAG+6Zusc6gHlU3y1q99SkMfWB23ni8pm4x1vIHDeV+bLAAnf+GzfbXBlCQs/00KGKhrL7azyvGR8RVPQw64upI6p1ZGeJqk+oEf5a7ouZGaHEwa3cxU4Flz1FaGu9MqNt2y7v+LzyRy4lAjeQ33DV8xWNwHz3hMa60fDNQfRCGEZt8/TRaxa0jqDSKl9K3AlhzfteJ/q3MXBsn7jiCw2hTFndjPvQHdix6+08hkA9TR1Lex23Zwo5lavtoOijgyolCRoHI6E5YsMtJY0u8DW2U3QmHwbubOc00tn7T1QduC+4ZTvmlA2bpvuYTYQ5/bDHnXcDt50ixjvdKEcmE4gxe8XGProy5V24pbelI/eftZGG29o251Ihvp3MA3c+sqgAbP9cM4IZwpmCNugmA+GWXZSee4ZYetp6bvaYzHJLvpZ9dQbNgNqObw5Vw9pqKThuLVBDvTdEXglOqHlA9FizF4Pc7VXFrHYkc61bghGfKQ/rHnpGHvYAijHdeleg6cU43j7vC1eWonHs6oMxSAyDGW6llxs32pEdDL4WAPL8RImmQrjDphBVURcWm2YM41oajzncUQU9zcY6cp11Jdmna0kpLLo158yciGs6bQ27YEZPwyhroQyYJOyVrC0Z4+kY9vFbagszrcrIdFKYDT1eP4nAB+lFdfY/cDfv5nFyvpCwOTR0iZGbTRB3oTzXfDYnaXrtbOEy7axC/ND6DE57Tj0ngWnPsgA8s58n7uMEemFZy9g1lvQw2B7QXxmnp210DFrzYOlocniA8r6WFSTkGdttwATQBnLG1mbMijRoQUc7kzbkrfDDdVfTjCT+Zm/+9JSPy8U9ytwLd63245oIr1MY7pnG9WpAx60XLo/oYUoa9qzaumdEg80KLMynm6v9flu032hRJoecRCc6qzi4O5D0dzjOrWg5fu4UnGHLkjtLcBk3bu1idUce5UC1i7YVeZcjxQvLin7h7oVdkMFLM5Tal2MjrtI3FlwpQmJJfbdwhw8vGANcH+wbDXvciKF7Ry0GHSiUqasddxQLt3gephtATyZQ529LarhA7TDqyygxvTHM61Uk5EIbMk+erAnQ74om1TZTIzdyI4bCwsiSovxJj9E7DXNPzWJTPZe51sM/I+iBeelvN1I/OMRnSSIcN+nHA3dXrO0cB/HUBLZw09c+cAf52I7xuvb7UshTK/yCEa0j5ST6gGKQuJTx+DR1Fu4+TVptWRbJCHro9DM+KxN44O5+dcALTkZxxvudfTT99kwjMExl4MaPHq8bLY6b+028WEjc6MygBTSH4U/cbeiN283cMUTL+/ZV0XT2rXuXGW33fj9w99m5XGW6dZy4c9FJlp0++6xbhVIkkN/gAikaiTMV0M30Rhkcw7Twe9xeGk9Gg0pfnheQEU3vb+lf+PWzXJoKsacVNXY3amGHpWbcCKxVmZY5zVcVsMIOKcioJUQLIYrxD9x0JkV71L4Z0tM0MmP5NC+iewtkj8tFK39tUTvuLlJTKbhS0W9ivegWnWc5fdEn3KQCUq5WUiwjPP1eWkjETU2+5sMCkK9HKJoUyYGFuxfM9fDDKTHcNAYr1nbwLsfNjALQxjt5XDPEZ1bVNuHBgA6FGblPqQ/cni0u3DyYaBzyi+xNafB1IH3HOKog6jiIGzOjLgyHPSF5+99T61jv6cy1R8EffIGMU9XtYmDs2Qfz5V0PYEdW4NPiHUDzwvI0Hk3DmJNLsdjvS3XWIvsz1TThaCjkU6yD1eV/1kIfHz6JXIthaZkJlYP4qn85IGY1nn6Ayk06WhkHluUwEagaxCwST3fRNPQyZsfdbdGJBfuKWpBnO3Z9k5zHomMnPntSmZs53hzynriV59nXs7bitMaYKpWz2bhz4bZ+hy7R8fJvZga5cF+tF2P9z8A9dUF9MTBqyMqsgCuWUbTSYb3r8TX0vK+PcgF9BXl8WcZv1wbLDffO9ufmuq5vIAL5d8eXYUspYQJ+lqWirVwDzIg7PWNGMZi5IoEUpcC6YZ0fFnkU6VrudFSM+hQ6l8ZqqEQaZLBWZdZ39tMU5d9wtzPJbvthkFGG2JlIJ3Is0vkUIR+1CDCKms5LdPsxI9pYJTmcDgu+FIJ9L8H8oWtQhlXGYtGaSuaC0UHOpqRifxtBF3L9Bg5t8YpbW7hh9SMvQgqK0cUIfr3xxTLR29bOiB8sCvbwCMjG7TqECgrMROgEstqmI3R+kxcDQ9OtEJHtpI5oLpUBhv6Jx8wE7sZt/XX2C82QXcOBF1YLZlF0Rjma73kVIIxhSxEYZCVzS82cYHu2C5nTmIJOqTIRX5wCxPmegubYyqOJAn4X2ZQyVv+B6FOxbCn0SeuaqbjOC5iv67OMN2ZfrowU2v1i7MRtTFPRSLhrShTLeaX8+OSlIkfLQ9EsbdiEbpuKOCvvlqVplegy5nDcDABpfe7hqfFEulKOn2dppEen5geVV7MesdrcEROcSSusxBVdFyMPNQykJ6GDH+sZaNHdsQ8t3aG2856B8HwT8DNOLu8jgJk1kh6oj7ELl16GAcOtMbtH/QygjzPAnHlhBmr4GACGYynZBBLzXT/GPkP8jfsOfEvIgK3Tb2K8wzlGbwAPmdfFXpaNwYBQOujTS+ZoLMqGKTKLce2dfexVRSvS5ot2nHFpx/4FzvbsgTueuJf3aAflwmvv7jtKmUGdKVSmowFukQdY0HuuL9AY+VihHA9lr7El0jZv9kEoLXrDLQOj0I3vmpqt/tmR9INKbRxVZpYd/XKoeytpQAqtR8MyF8pTuIGIz9k+btxxvek0fB4AQ+RawMcgd/exCloTwZoJYDrH/hkcs3knttJB9/S+Pgn4UQOaxWjh8aa2PdU1KrMrWj3YNO7i2OX1POh+d1gB1EY14v5YQEiJaOJO+D6dLxc+MaUfip9Z29fNQO4+x2CUFn31oKdVPJoPGGdMABhp0KgZX5yqtIJhpgycawnG+xtsfNdRFDIEnxamIKQALDa5sK6u6jduLpZqYwYZbHP0555PO9SksXZ2QuVpI+2imle/1T58DcWlrmiE4bjL6EPGv3APp7txf+HnleT9D8KKaUepadgXbK09MlA7lUshq+3BR1NyiNyJm8Na1g60Avby7ytjgussjOcu76KVhF5c+dvB6mSYJ8IeVtzmSMwwt6w3bh8+ZNvUmMkg7rrnYlFXK32r+FzFzx5Go3G7rfITIRvrelPn04e9l+7tn8zmys607Nwc/XXhq2mb6AU/qtSq0GEPxYVbK8M6W5B3BQtN2emWbSd2o00ySAytw2iq2OhTf7B5cDmqmsXxJeJH4HNML6YU826uIL2u4knXSYg7H7jPcxf2cO0cdyZFOpfwWKFqO071PDMmppLF3/7+qFQ7FYhPjptT1+JP9pp+KYX4+1f8vYTbncztvCQ99x/8RCoqrBZhUWkTmv2iId5yNnaUnGUi7OsNd2cjlANx54l6NvvgwxTQAbP1zIPb9KCPvnPclpOUzDSrp+j7B51Mhf6kvbksANz517g15Jzrb85qV99hS49X+EkOa12j0EsbMh7qybalLtRCDqeH/76uw5wfh/h+7f7DF9eVIIk+hipDVzpnQA6Pb6BS2l6cUsZQ3imQtiiRjqMa4FDGNoVFXNrKEKVA0yHRqZAUWxNRfSjCcjVidGEMHHbIQKohL+xmNG4GLH9bNzismri7YFVpIQ1c41MqJqvkH1OS3iZ/+quIBovg1AcZAce85qRBmS3cxZObuEedomQzzrssHto4ujO3qMhsRkrcEb17NI/Tvhbu7hO2NLzTbhmF0xYBr3dofC5n04W/OXQ9vLx1/kPzuzxbwydG6XmOAHNwU8chrdR3PCuz2uzl/if76uAVtV+n5c1p2F6gBjkIRX5KOLsW5LjpXB131xfpQB03HTB1iTgIb9pqfD74gjWL5V34oLwnjQLASdW6mKOfsDqERdOOcA4k6xCPS0/2Qp022OT95i09IqOGKlL4oCEbkkqVmXUgXKFMiTAZFuJD39crTl9w1+a1/OtNPBP3IAqqNgv3HIf7FGhnP+XIta4iEcLdbZzraPq8FrH9gDke4dYQkEVIS70zVeNhVnAykHMsXfKaoA6GiiYt5tPogkPPswuhF4fZ8CU+Rw8jx5Rns5a1mzIowz3X8PQwRGXiODhVKzC5M+M9sWStCZGev+Befcow5QvJwwAPXaJTiSrCtw0Qpw+5CbszDA2hSufl0IgTDEDMIDbuORzkc9+4egrFIwW1qj1TNV53jPMp7SPfe99DgIcqKnsZuVIsyPMHUkur5dmkpFweTq9bKeJtKyUrK+lFLViG4Om34WbqVbgVERUlCeUdtyKJcJsDYsNS7k5FlQEA4HmjI9UERqRs5wVoE9FweKV8CXMcLqCO0r16k9laoA99M9yZOONZW8Sm5IS0MrsZnTVW4SYNpkM3KhO1IFCdBH9a1jv2LCGrefIEw2Ee1fPnz3O9faGdyNS3xgT9t9ojbmUqwJhp88DrmVnZQK+ERmMGek+ImjA7QDuRQ2bj3utver0EMI/ZO31fYfjdmcjO+kxe82r4+vJSVWuvD3z//8HbaRGZmjeLZ+2JuGW2Dw4tRyOF8/TNprpGlGDYcwFzDwDl4J6abzpvI2z28N5WvHYUFACFztPCzFDxZwKLwv2n+0dKX7UHLp3eiu8U9bLbznCYAckgGcVWIbfbuHRvT4eWE7qmspPGzsIYuatvDQmYeTXuLP7eDIielpiz60VL9v2Ls6LFeUpvrKkr63xSi5LB4xdRDjPCcPcM3qEd0JmshltZxkVGsx5iuLl3yAu+JkcOSR/yjnLwjim6jw4GvoLYcbPg6brZw7Qn7lOQv2/OiJSOI4YMPHtlVtR7YG4FKlmKLZMAgG9EnO0vYvJOz2Mt3e6x9mUd1oXCFQ3Yx6rKUthHCfE2ppQj8KFMVOTrtK6VKOFCuJRWhQsPsFcAoirl22ihSJNIYQ5ctmS9XN/1LTJvw9UO6DxntD4cQynP/Vy5ymFOr0cx5TrEG5taVj2z5BGtnh8ZQV9HpZwdlftk6JOBNW4A+Hz+C73NvrOyzsIgvpIvjbv14P7zzWMp3vFEberGLOZZ2wxKhds40rQxU3XcrI8Jtw37hJsrZRv3dX01ddvLvQMXPsIgx6e+73U/cN9ZejkdgGcaAM/EbV3q/3Y23LgLW9bsljJ00ytlWjzrtnFf138Vn6yEUH1d1+fsWym9/SIzfINYR4oWJCNmR9UjkA52dtbgcDyhSjoE2IQKjPYUtcA1CWhPaArZ412LJkcL2lQr1WqBJDL/zvLhALTGQbgh3BrDanaIhasupgZSs0K9twb2LA2fWMtfcwx9L8fMFJX7Ty4rUInR07l4NsB3xz5xH5yX1LQWc1nKS2cY5K7pw8CtyNyp7lX1BcrssMuDTepnIoHaINfOghhqSt7XDEjk5QDWPprMv5P1MOPTdCf1SiV3tUk9PsPdfxr3yjq4CTCqX31Xw9hjZDbrtHEzokfiHLFQQ0xmOoLmGXM5k5VtSHfI5ZGhQBmX7NOGimP3bgXrHuYHzmzNLWc8cR8HQzv7xnWZF6X3gkhjNFCF+wo1dlfx5URannmQJtwbXrk+c9mekdTaBXr2Aqe9C9FOgGB7h2QLXcYkelOKwmdgDEWmlJ1FpDNmJguijOVqTJfNvFSU0dw8R/oW/egYNI9Ox1cCOXddGPty5CA6ixmOzLK6phXClAFEtmKNbcnVovZaMNqEOGW4OQyFUtMDpwxdh89wCq54owQpy6BO5JVT02sjovUCxRd9V/y0mZ520LOwzvsTqCXJnSEpYFCTL+qU6fRwxOioWt/RufSiLhhu6jhrXXfp79FPOr4WZAXE4JoLZotNgEd2X5k89q4UbhZ884G7s5nkqxH4fDIo3+3MUPLUsPIz7Ji4//6Q38xMFTHjpB3ByD4AUUOpEM34c8u519+KwFSZStcZCNPNq6YZLdIerao2zXMzE81bB+A0HZeY1TMINSanIap4UwxELwIK26Tlr56zTtqgTNByCy6LaCNt3ORRKrWPi9O9f013TtyHZovoxZfHXoKdeflYdykBTCHb2CpAxOFLJwWdjiubY5+g8TqXih+gojObcoOrrdzZ79M85bDSC5MVa1A0InJhyMUy2tMu9QzIZNpOZ0jn1nziUK/XxdzwTDbUT6f9LAhHkEYarNzLwMFhOYdZ/TCDl8u7p4RTDi+NEpvSzDldS1mf4PfRe2CgoXLbE4cjvYbGRhfdvNEf8c28S/qdcnqgLk0zrxUSPqNaR8BLIY9TMOFCkse80GPvFMiOGne9XLkUP9vZyBPbOFasXecZuqKk94dsJxNzindEWcus6BF8X4hHfkQg7hRffKbFI8VYQ8GkSCdBoRZMwZbmAvPsglQkPDTcP3BjYeMDXUBzGQ5vR1wMGhFjR+rALSPNdqBjR/HGbTp2cRm3RVI//tBqLb0JreSgsygaF/uPGmuPgqRFag0biV3OgLqJZbgs+jXvlE3IqYR+dzytK70oTdms1cgaV2GXI+9I1PteaAukqTYtVm1FTg+dHbiMINl1P8ymBm63r4j8fq6vQvd5yaqnb/R2GMC72sxUrQXWymHVVr4RKS4gbvRiEVM+MhwdjZEBP5RFQ7FkATLNtWV5WpTS9PkKuAKX3sJV94d706MgSudkxYY9MXYpCrdqL1wjULjsgFlV6JX5dJp3gXwwJc1O03tPQ+OWw6Mjt3MXVLQrkXAoMHGn0dWybdwt6oDh9o1g5cR1sli0DKSk1wcni6SRGV1yaOeoOg2fBu4eKsnBiq6ow4s/K9Acui4VLOu/0XULxKeyAuoJHRF5weUBlP+a5Um+V6Yz2jPTx8zrAlDZc6X4nB3pGlU7VM7wJPv3jI+6Eq2HnGgYhenSyPM2ucpw4uihD3uiswDRRNzUaemmHWQUQHypq2Nn3chBKt7KuLPfQhY4RT5GF4+oOuiW1FQUlCNCC5+MAIVu0dIVmRL1/wadC696kY+PZNV4ZuEsEF2klMc2mo5Wt7LdjJwbN9N4tLE47rylDB0tBLxoNidIvYRFVEM9C6rdjhIO4o4U3zpjIkuoQIyczS8pFI2UzohDAsdNHaHTDOC5SOzw/mQTvaaDjlfStexGDtEc17nfipT31XhEx8Ith0Om1hSp2ryXjju32ha6RkDcdEDMIJo3XLF5fOctPhzcnDGE+moHnY3bJJ6466DmPzkjHuuvQEYusvhJmijLN1uSvJ3JtG0f/gJ33vFl9L04nuT5As2ujm4VsfwI9FD0ZSZhFX4d7gJ9lxZdOxh58c42OJkyAcejdlGxGF/ZgU8lscqLJUQVKqnYxF1pa+NOixz1NzMQRejy5rbasKvylpGUYfmb2M2sKRoAhUHRmovPDn8u409cX2UurLC70mosXLQO53tCJq74WLq6cKOHDAdTB4DO/vhqS/KjlZcO7PCU05J13SIsnWfXg6DpumPXPHi4M5VbMzeXxtrCYTwTbjoenRf66WCiO8mBsOe81pHlNy6M10UIB7PN1uejux/DVnmC29HQFc4gkqjWUy/4S8dwP4vV52bR00M0dFGa2YRAVHZltpeG+yTmgYwrOzxpXM5Gzu9XgdBSaypIZQo0XI6lPKX1aTzY2H6k0cwMwDFWmXe2sROYn2Ak1xyhIqkUNdS02j/89wJXF+ya0Y2DR8MJoznfue34HripQCWhfu4K3etZhfPiUOG4Q0pKGuSwLptlYP/Kzsjvit50sJbtjN8lb8ediqiKemZgjcVx2zQy2xVuYAiHQ0Q0D3ymgjgm7iPD87Js4gg1GbxPWc1nxOius6B/Sk6BO//ArIT9+u/igbWTRVPX4hpn4zaFzNk26VImHEbvbGeTAAAgAElEQVReoLB6G2UzDDh1oy/Quwy3HjWbhvplXfCvzOB+4DZ7ztoVYtNIGnNCQeooo0VVEsLpzrEu43wuE3jE2al6WUbCirjaAiwNb4WRJyR9Sl9p5DVGrFoIjZ/pp1eLzzj3n5rq9QyonWBYH+0EotsWr+7G7VGq0uQrvogI3MktyCwN2apKRQATqMahFVVszQqFrbedI7RmhN83bmsDifu+z9Z2kwnn5OdqwyjcAHSGaF27Fm5Xuurv+nwPn7NfrP3AfTgEBQo7QZzGeFXRTpma4FudLNtp+/QwDHdnHpA8VcuSnvdxCACGnnZA4dmlnYNppWcmPh++x4ZF/Td5Qz5jegUG4JJLORm+WOi0R/ub2Vz7vOIHn1fm0hhYPO61JAy8jrv1GEE7PXb0RUSvewiABR8v+nW94CBoYQEyXLByzls7SmgpMtNgeUMbx9OJ7KPOusAygWr1Y79M5hipFwBP1PDC3HV9i8lXp+ZHvcHiroSgOg7EUJSSHogsVpqQ4jorBJkFoRhOLTEFO89m4TdjN9xna3VPQ2qjj22VJi1dcGU7jpsFsZyREND6j8ZtHCe9A7cvFe6ZFw8EA/dyKGz7DDeI08MQtFWe51LM2aEOXG4cpCOMlqjhFjRr5HUrn0J2KlK80NAZLNrn4B1xN+/jX3AfJ5lr7wUDRTAo2TBZegwvMDtuOo7ekqDgGgHui2lZWZAcAZlZXOPmdcSFuCK+EfKBilRSIjauhR3AWWXY3ruVJIewD3wbj5KoqxU0uemKXjMZhzwCdUWZbtaBwwyWWY4i9ki/Qs6twHbGEXPaNOTMTH8A9fHATSNEgOsUzm+dAWnRF9qj91Qe6ypWXQfgB/DoHg1DqsoOGqa9AEgOfuKmD+j2L1Nsx01Hz37Rf4sZsx6FChRyLDSW6zhrL9xxrH19qAMLd7RRMyhp3QZne5CVORRdg5YpH77PVou1Lo+u/qhltdQlyRftgPQCLDoE7/fYxnWdWRo/x+SKU6TsE73CcEcH1sAMvOjsvHmScgjnc9vvLaMO1pUp8FvP1JXkFG7czeuSbaatOw1vtCIDHxbDvJDTOnIWgFQR1CNjoF2FphWZ8qa3yeQy1C/7ua7PiFKXVXoP+vMUr0cpGyor8rZc6E7XWYh2nR2jiHaO/j2LSyYOTu9pmo/8oBJVW6rIj0zMBMSfEeLTVduVo+i4tNI2B54+W+OSQ+IKwom7ea9UnhuPHri9fmD7UNPl0zIX7vDIF4Z79ku+6plX3Kgo1/WglqdpCvkvvPwekzY9bxnAwi2pKIkJ6MyW0deStxXhx9/aRUz54gS3BHznb8RVQ4C73qtlGxdBm6r9P9Rr6XvpvuiE6Rr1lPZysCu7C9pCGObWYel4nVDHs8DM0/7JY935z2Fvnsru0Te+nflGp9S98k4KZM4FcWu40UuFK5ar6Mjq+9XPXt8yVi7HDt3r4iRSn3e+amZHMyHihocSj1osRuXAjTLCuxa79NRbzjZ82TyfCx4JZ7g9OsGU2d5jecW3olJFWWUI98DerAiTYR3JhpcoBEb9nuI7M0Tn+Tv/kRH3u49tkRTH+/7W9eEwHDdxOk/CyGdUNtzX1xLWWl+j7IefR+FNJ4yB8tYCQxg/Uv2N7BNdg1Fxb9UmgDAaiGMGLUXuu+2np3Ibd2dIjOxXTdCZARvdjrp5XrZiJ8ppmFpFyiu6yDnw8fn8s2tX4zbnfEz2T21cXhBzMc7ikS1wQvZuSRoCvVCNi33fgS8jZWGws5ZU+4qIFhWOLG59zzZoZnIswFAoOT3wfRu3RdsQPcJTBtWZT+MGC0dpPBGGow/MfuTVIw6TGSWE25yUImFlDTSe1g5NIYt29mnpZ6/Ug2jjMyBuRiq2mbA0+FafijDOG47ZlSJ39PpcX4tkjKzHEBkFxVegM5iiwflG+hjNGnfzmREuNESgbTV/OZtzXd92OIVNMmwrsghKXLcwpeReQ6zCcXBHR3DiV+ZNWV4Ld0gnW8eaRyNzsoykf28+S5do4KU01/XRgdYt12JuUvcAl7nr9Ak6d+MxvftqnrbAX5+zAmwYHxhpyniuJo6fLEGcAt/NwDEVj09xDG8RnnPokLKcqMd59/k9yWdm0E5DxAQ3gdETs3uLwhbtr89HuOlxVcuIs2nuqjoIKxzIrJOT/kSz9w8Jtw17vAl74K7s7YHbtnQXTs4YnGv2ZirHfdKVxp2VSWDOOF3Xf7VMJDLiJw1Mi28tVUaE5NEy5u8dbwfuZgWuzwfjFKiKiGdPw8mg7r9/GjdMh67r7KId0+vNm17lOtVQQe9qp9IaTtoDYe1Qnmdm6wTJm8ZkGfaQAUr0MXk9Z9+g75SbVH8t7+KlCuhs425QCAPZp5R1ZnWc7HGgNa2clmnx+XbZnQUJ96Hw2+M/x3HbGYIFpq4fBbtwazaCymVTROIZiTnRJDkXZJ5d9992oCpTSwDcXMUKuxddDqNWAcqHGGA28m3FIl2WQup6pHArgwSAOnn64O4NR1F8aOdGljFqh9aADLyjHsLhTRfsGOGOPG5cOk28PuSRTW3SwGlUlxzLmk6jkMdQkY4n7F0flxbByYmSzusCbp4y3tV7p8+nAI0B6ppbyHlqE9UvkkMYe3WlUo7OlnoTWHR0B6fsuRCtN28p2gdk5K7j/Qxxf0tUPfQ7DryCRv5TcKKDB3GPYRMhWOalnAFnyKDCdpZRt1ORMwWaV3HBV82eLK3auBPxuXD/+WI7SMZdXO+6HJ3VKTp/5aCEOy78AfnFGIB2AQ2ZY9OUUMvTFBTpf7ZcmYbTqOI6px1bG772QVOqxx2f9sjg+EixfJxKhQGjqBS2I9A8YQqitesmjMY0GhtuuQHQ4xO3KfRxEk0fcalWYtNow+OD3SRQB7XeY3qwBSYDVx+H5jmmLSiqAVEZ6KxiRLkRTcsxnIYsCGhxT1LaZXhHT26TC52ozIfTgxaBKYpb8v4D8Hk4cmVOP3GbTCnYV9yc/ehrHTZLDxX0+oR1LWJr1OZwCmtF5PN8rexMWNDsTIO6cMue7orYFBpn8lo2WschO7AFjtJNBgnDzawoejs8+SLHQ7o9GSh58+8pEyAi4usRmEY3pvZ8XM8CXzH7QqdmWpZ7lTergt8o5sihpLIEptzsF3XdpxXj0wes4IimHQby0GQbkJLvP4gSKKf56GzsZbFtdD2fPpQECWRnM3IoYESe7xfRYiO1AyhVFe4e3ngx7qSJrQz+zhVG9LNE3ZXAsrvPp+4rfnJ5NnHX2Fv+M+kEvGDY/zUA6KECXnH7bM2J0vWwRe5ecFrBqAi5iJNOIllsPzoXLm8fOjBLsHY59XgMyQqYVkht3JaRJeU0GNR9MhoHC4nnVuGmQzR+Sa7B5QIWGKNmN0yOjnvMOhoNpSjwT9N49O7g/lMA9+EgqxDDkRhuBmnW+o76XPiLOGdwdgoLNeJLe9376HOfcyVOQZM5Q2cNNM6Li7wKtJuhVPOex6y1N4cpG71u05a2Zv/8Xamm+iqpJjDTw07hj9DNUTp1xCGlR0XQTtuPcdIJdWrMrOLQwhWck4uN2/lhxq+xMaNBKbk5iH6yIn4YD4lbS+lZh/jr7SNFp1UszGn2Nb7/48CrlLWcF43Ra02n7VnRpziYSenC/9fXlS5J0uREV2QtD8aL70NhGGu20yl+SH5E9UBj8A3dVZmh23VExCr0hWJI98qBNA7drg+JY9STXv6krghF7EasAlpXPnQ+xXIQoIhDkWXQpHNSHdWItDY6JEPaVrAMutOZbtDtCCyXndABStaBkIiEA3lTrxNFjNzMz2s9f6Wbmca8lddH2fNuBDPKa3BqUxGRtGqaE/K612Sg0prnHi3mvQk1p/Y4SrmoqHWhfJlNRcEyCpHvFgKV0sCGfrXYFonMUXBcQqReAXwV5RDPcBCjSesErbyQho6PlyNj4WhGN8K+ezCsYepLzlU8PjUOadfIEW7KjVGU4+XQMwdt5Qi+kM7+O+nW+qOb0F+3zM+x9R4eKzFl9WThfcFGP+9uVOUOyjud4lole3wpdE/64xvEXoGCc27+zjq9CZIF4nTwpvv9pbfSg5Apjutf2igmvsRGzPrSlI3Q73dqqWDlzxeggCCDXvnWeYDXTq47tvt36PhV7zHd54QN6zuUTaDLdCR1cM7Tn6HhmMDaHm6VDjwpP01HfNWVNljkaj+uQWsn4joK7g6V4RSJCvjoFSvqYCP/KC4dguGzIuEeJVbyaLs+QlQxcIyZRnH9tOlWCgXTlM9VLfvrBG6hkv2dDS8LtHxOqEnSrWGHv9OdaEzDTXs7mpRg0wfPiJTW4ENqRfiuh4ctW9480+Kiu5yrk293sACwN7gpEpJuGdRGScFx0t2/6LYsgy+i+8uo9+9XGkEunzjoRml2zMmkDm9dRkhKgaUtK9FdX45Cq97V9LX3iDp582e/sXqTDutcTnfT3ahfZMGZgWjW6trNpP1RTsBt31yt6jJ2Y/UxYcy3dsjjtTAGQe3AlPKyNOI930HboIf5KNpOdErI3F2cnIvOPYAcC5V+guzjZ5cFY8g7Sq0DO8bl7iszL88OQa9Di3fSuPfdb1uorC8kDFWL9XXel/k98v92g1cLXBFOkKVWiFTaRQVX+rSKFxEB4QwB+Jl0cstb+TJFfhewnXKV6Vqklp0hRmGuTxDXwv6VNpCP057erz7saAwqedv1IvPCaHP45V3OheHz0P3j7+z7yJMALbumN+zcsicPxqD5nOBz7ZWEy4Wr+KwUJ2o2q+forbnxOY9HAZDB4ws9sd6UQ2kKEouWzHtye23gOjkt6d4SA48OuFKm5ZtcKp3opKDoxsc7DkufPco1zfzif9MbS3v2YxwfDuPylW9sCzqvDtcJF5EJfBmN4UitAmBuBoLWUaARGMZScHJVzA3fQDKpaJLZ+vsGqpwe2SikTchWqfcTHIkQ6807GUYH+vb9PETkbsgxEsJm/FExDIyA+x3+DpbbLzRWCJooa8uF/peRmSo5G0/jWVTV/QwLY+N4V3ERKCsUpgDg/dEVkFl0U6q0OrG/VOTWXAjp5ne+6NaPIr+Lh8OL26hK+hC8Ike6QQd7031m1ykdZYWepL28lCfWUflSZKfhMwsx209Il1v1HXTYDnNmifKHgmGifacaMZEa9kY79e/Ixt57Q7ipixfTyG72C4kYlhENqLV6zgGvXqOH51mSi/C2+Oct0rfhGRqm4nGxZvjtAKxUJRSD/Lty1WV8OYrMv881QKa6QZXX1LGmXber3A98YlHSHQhkUzmiT1ajdwGXwLxVO+hqft+eXrTVzikkX+qbbhe3JBsZLnyoK6AR9Oz4cHiNA1Sjm4GM0sfymTytmz9pcMU6xSg1Tu04/zoCzhgs6kr0xhvORQ8f/1d5O/KrngVgCtt98fZeV8g7BwFRqCdSTb076K66T4GP9WG/bzuqvb+EtB6tnagh63sqIFfKhUN3BaLnS4/Zkez3ovvSibyWANBz1eZt4Dwf/PxhNwRTsKraA0BQcC7aUmLFESrdCUUbLZFyuIq834oK9ryzuRaAECo8OVeaMC0NtUCPu4J5/wR+gM/cLMwzIoI0mQ+Y7r2ns5bhjXcd3DBQ7a+a/rjqPLsOvrojspsna87l4p/qH4LKSft42BIvqdRL2xfd1t7ZE6BoI8EYCbAIWBw60sHKS7dSENqy6xtar97FyA85s2wLm6agG3U/R2jVpDNAuMXNz8UF1XEvCHmyCx1arkBLw/Ev+32VHiiaMhC2T35/6uhMkkZ7PUyD/0L3dQ0lIPk5VZmgnINRjCZGx5BTz9qUisrbqeBoN87Z+hJA98l/VX2kx5pc5mujsJt0n7Dl/Z/+vO8ftQNfKi1KzJPDSI+1xMoZZIFQjgLydoSYqsBvVd/CaTNtvR1dUMcz6HU9brvRtvtSvl0xCMW+N2DROSiK77b7mR7MEeJGc/yXEr3gbIZVO7IMP389zKeIPqzThpgAT1pnP4HvmTISaxqEoGUDJMWsycgodz3hFAfGwk5Li6GzjDWJtlXy8wybi3qwst61TT7+NRAV0bNJAeUPiKfd79SJkm7x1SmmHBDTSi5afHEnCeWWdyfTu0I2LbidHTSq5CCNldkicWna8pkdNZxXaCxlK1UpcsA/IwNoHKEBtdaZFlBv7HCnGbFRFFl8HZltjQzlQTilMLi/v4gt6ZYi7GldH1euKSxIaRyRy4KX1/MhHvLcsKeybRi+2yPbm5YWaWhYgJjky39caHz28FIPfYXTCWbTqdUW1rjVfDwoDX0rwwEvCUuNCFj9Hg/O2X1GEkbhKycMB3FFNPIgo0LSDULIR0M6fN5Ft/hklME1nR1vn4N+oLZuv47oLoi6kmK6celEfn4Knq8H4vbzZ528nAsRXdYN9uekIUu76KBINwfuWvWAXcgiwt9003lcJ7hRZ8vfpcMRKhDdlFfOBtFYx3BO8YzQsrxOGDHlKgdHnUI47vzDyv5woO4IeZ7nYyed75ONBd3Y1nhjdSTOI63SzfLSzeW+RgZCzyg/8XDuX2E35LdX9SYrPjCsiQsoVnlX8cJh8HCWbG1lW02RJ1o7w5QkCFZWwn729BEH9644SIu+RwZQWbi2/Xx2FC66BUnjflRQrXyyWNJth3OjrSkyuSPBTUBq38GzDAqOQTfhro7Eg6G4KNe8RoFj9ny32JH3nTAiFCnD9N/T2V7Ig2hoDVk1ruPnKu1gahJKLUl16JJnGUJqMPLCKGm0K1vtPCxPHo2co18ddqSiPeqmO65MEOXZhdPtcJtWNPXiXM7AqM3OJX8GfYSjDf4k3Zcj5btWN/wuXvzln3M+RlvdexZxTJkGx4H2nS9CJifk6nQ97xU+dEDel9QH2HMTDx8GOjKcsgG+7w84eVcFPOeB2yssEnYUhAxnGMFQ4/VYHZdxaz3vCjtzejJxDs+dv+8uTTIj10CGFB2PkcdkQlvwqtn5mAVSLM3eMr4HFTNPLDpR01JLt7sg0HrmTIn97HvTTfQEfgY7dLP84rKSbmyL0PDb0fEsvWrLgkhl6T/Hsns8iSl5n7OFwFnrGM3SdA50FujSIpkE3fy3OxQjKw3IgQVKyho2zpT7IgryEL/eAfTuoJ0ReYinWJr5+RnHxkX3reNLd9XUvZhC77Olo/1K3veaFsqHvBs//ruu+8SilNiDUwi66cTbfBW6gWyhqSfU8xO6tHytqjXy0YeTdK8zVg2nMHRrmnhb3AIRPO8D9TnnKUGbjbbOh7bYc55r9yEA/Pz8G4zOw4z1/FEsIXDynoKze0bs8YloVBPZqOf5+HUJ3Xs4imc2GDkd0IleGB1huKb8igiChSjofd0v3ohO5/D8xtZ7m3Rrt6k3UVmZGf0ij9Q63lgPtEY9v+Ng4+XT+fxjnE1T3qS7L7rxRbfpXceaqcJ+DltPeHd35hjgIxqmKPdj1xzH4HHHLdfkCDtRlelA1gpUZFOAKOnAERq96RYvxTPTzTkYpZecxylG9oi2rOXEwbVdSTcHmhv97t8u/ds9NzE5q9Z1rO15PiC7Fd/7DbmQRwh+OwhYzynrfTb1ddMDTmnyGRrRLmC6eby3NGektpnws3MjtZ9bnjca/fNH6xunetANfLKai6q55fqvKchGnz5SYlQJKhIO0ZslQvBobq9gWFcgKqiNgCXvJ0aRtcrv4bUBGryyEOYPL0/XYlHV+YaeT29fSfd6Hk6ocv0vC53aol7XwEz++HvOu+fB4bgcMiLqNAzf6dQKHqteTYHpueY5ku4Ergwruw5C5Mnnf5TG8L+cPzjno9Pdf+XpEb0vuhWNvW4gHCm7NKlza0iiu2669RKlBaXfDXLbEfDH7fvUDXyl2JJLOLVBxOOwzzl46XhfrplOQQ+Uvt3zEt6RLEe6BU0jnhPfXae/dBZOPD+d/zg9FV1Bx/sG3aXnAFCdwrbDNQxvn/PZFuna5PNoYpfBS3pUwAfd7ZyZCxmlfOWp18vpfkYONLV2qakFQ0atxIg4xgZDeMXzAXwEm4pTaDEcsIL4d5U2r8gAMOoQ6pcjk9jPIlzruxLM0t3vGlJc8qMOECF+QQNg156EMOL7sJ5dmw5eyQjr6j8n7SzzcLxrJM7bmb5I90x3OrEmv9aQFpnsF/yxpkMgL7eAnWd4lB0kDcRrnXd/H1Lk1qW3QNtR1rUGPkXOk9AxFXcj5UUCecw9SPu9RG1Sv0BBqilpDVHziPQgUz8dmV+3bI2gg5aQR9bYzBsf3UCbSdldbilQKXWplo833VF3AuCLkYJu6gKD1vt6N2szHV4xTVrZH1RGoVxa6cG3sh/NjZvJ6dWchoBIITweU4sZITXC0DxFCE6blbjGPcuT7ykaMz1Hlbc7gxHGA0RXVL5+l2QzLEFevcGDR+zRVRPpwh0hW89JNMMo80Yd5qIbUGrEcV1Wu+dvhZx+bbQUQkW4lRudtERauWbyKlSXfNoPqxIu2S9PLvWgcifd4eSKRyHSqNfRyNna27PN6LZfODDg6z3QsFZu4Rereap2T1eC2xBEgCPMPJnpqAYP92+Sd6F4HaLQDHXEju/ujtlYL76Tn+13V7eQjunm1Ot2KnIMhWmXxLXyjo7fObyn53vsO4JtFOlFR8SggnV0GhdVH1yVdUYgF5Q8zbdffn/0NPPgSBn44hT4Vblfl8WCEurcV9h3698iYkeCSY86OFr1KmcYQ04Zik1S6L68LKgQgYrC/4ARgMLhaxQJ5hM7tuw1NaAU7VRpXLvfH+A8OpfCivXu78YJvl+XLVs28HuqhMbM4xN0ByoJuGsJLd29MFULJ59+9GghtqwBkGO6LxSBjJy6DT1/VAdSMBHdbsW/Skdqx+3Nk1I036IrLFO3POumm4i105FuHepFpG3sbPWcmxkI4Tk+Fc1rH7mbbyW/6tDcG7RdV4H4/m4XahGcOoQFnlrf290q6u75CkJkitBGzFm8P+NElI54d7dTJ9rbkSwyTXo2RTvn9AeoupyBLGQXEAroz4HmYcVNOLb/5TVq2TueaNDonygoEfrWHJBCZ6OCFXpHgu8bzTyJ1kjFy7WqbUoDCG+f9JjuLQT9opszJ8vGttMq8BCghb4L51hsY4FzDgvykW3k+dBNpDFKO4LlASbRkgZPwe7fdFP473dHyXRDz084WlLkDkM3SDKsuOopG7np/BVdn48mLFFnDWLfGV7Y8zjKpIUyiAyYJphu106w6Sf1TyntqdiYNsawx1J90X2kG01nt2sJiwfAU65spEw7rnmH5zP6djgVzWBg3dMogVw14FYmrw/cdvPq3ZzU7Za40dGLruOb0jnsGM/eSUutkTrzq3Y2n1Ig4OdimG1vUY8LStheY9V0WnJOR2Q4NIxdgKLkmRrFCQ8nGIkeNAHAM+/hJYWt+L8OcFALjJDtQ1XAPexS+n721cdxfjOnxXwVkNZRnOPo7DSMH49awwphDpC9W2Uptotu8oR0I3+IbPbblTIp1DoKoiljxhgcU2sNutDHPF7jgR1rDiHN/oeOtWUniWuyk1TJbH+nYbekuwp5qbIcxUU2c+aYswilztmO+fG8zIg7jkNA49HBPEQjCLotb3UEKoLB/0U3ho6zt4o10Szs2Ob/jYOIiTREd4VeJN3WibmIuHTE3/v+UdrANuv8+5tuqFjLdEeBcL9A/il4x1Qt13B19IRsG59C4Tz/uAaXgISbsyjDE3rruyKf+dk9FebIIOEKoiEEQgUwJLcwCZE2ulY8B7CfWMjJNblAGSlHoBgrRPLmgc5TFDyvjSbzMqcF5c+cAoe4EtncRsa1siC7Gswt5Bulwe8z6kWFHQgE0uG4wsDVUWlsR2DhK/PdCp5QhkRtDXAUnxH/F92UETEgnUeMOMt50Wuits25AutSZHdqe5lRjPXPmvjV0RF+yoZMAzEcX+f8ku5McWmYj1VIdGO28QulcmgNw1tkVwcKkHIoiy7VDreCGtVi07MCetMzfp5tbFTFtS3mZSIEohXrW8i1RibFwiscqLLj+b5Gi7OuDlTkFvznnNPnnKtIaMia3p3KcxegnFPjWrSUQsZ5tzDnVKfGnVo0WLmdd/4IejpXnG8PY+/ZBRkf4feuyeBlDVYQ2C1BCuSm2zkeFa9RosO0QL9rCoQTfKKb9RwW6bbOsHB2V7gkTBvQE3Ut0rRfoADXiQBNwRKyK1dNuo/WLQW5nPau8/F1kZeh0CBrMIVrW+b9Ne1blo/WFUYEdn7C6fpKw6S7FRUlV0bEL6d8eF5EIGU8pB2WN6NposfHMH/8/xNBxOg1U0CZWNJ9NmC+q6v4vnrA3/9uvQsJCMXT4XjyV3Q3xKfniSnedYbn+cfQxXrLId2tZVSVrggwbx89JovtB0C9P3+0gMkXXxO05AJToGKlt6R4bKnZu1fNXHuxjFuO+GYWhBjokBGpAy9iydzbBTYOS0F5aoeRaGfl5TT2fwVbPW3a7w/6fXV/x7dSzF6QRUsIR9OetCQvHl5AnHTLwTESb0GYqtZ9wcKq2gKbC6DiCR3bHmCSdYw0EI9hw99Zo3v32oX3549kLs/Cz2E/F3MsnIaEEAKd8dm12e+CbrMZCr91hbJ7VykfPxv4ojvmU+jEXs5EkO53neAPeMOa08dG94948v78W3KnvAV4uKYTRhe36GVg5LBiABXzMZyYEGzQTWBwTYmK7mMj5jPp1C+6A6nkjIrQ/+g0URnpRjhvrXrR3UxtQzKZhQ59H2Ww2dvlAt4XeDzxRsj28/NHUMaTZkQK6/nirItXg16DSgbq/LmIM7FjYG+P4edx866Z5MWzLScwJxltAUkRkGsD0pgoAFXeEyq+7549sDSs19bWYeaF2ZqqrcC/VvIGJ+usZJ72tCIn3UPrIyOyY/q5FJfph6OjC4ZXxZ37AlAyZO6YVJq4uk5kx+sicw5mPptTku9F59RRlo/lWZJxsj8b2bjnAfqcHWIGjy0ArvPAOkoGNEVfJN15Bpg5PQsAAANpSURBVMfrdxfpzvmPe5iO62G3BnCxNIusGhvgM1UIj9SWdJ+zk5DkcxTUVQ9LffTn5meK3ANY2uuUvgFXYTSdSYxyz1d4idXJgiUILF0LGh4NmvTGwbP1og8vzxmnvQWvs8aHLbZsROOLOM6KKhkHhSCXSWXtFY6q4x1K3xcTxTAZeYdXZ7QY4enuUWBzzQMOXM28v++juLaJa3k2LHnzI3A8nv2J3YtVvpKgCngXF0jAHfQxQ9x5kpil0EGqC4krDSMciKMKeTtOJ+mmA2xk5whCP/M9txSpzGeNUB0rorvN7Z8Pa1DvJadbDqa7rJXgHhJt8IqpSDp91jX+Nsz2m5+1EZJHCjTmagZ+xvpWy6d0MnI+pat85lenrmsMTx2cz3+EgXzTPTWga2ZDf7Mhau/HG/aADAbWcSNNcSGeu0XUdz+/Ka0RVkmPJnBvuvt8vthXOuC3EBsS9e4CMr2r5/da1nl8qJyuS8xCvBWaMD8iMn+EKowo5BgSEveXQwmYbEa5jQZFKkLI7apowiyfl60uRzc5KbX2WK0uMY60WAnd4789sJWC7/dPOLGoPSRdANT9UUQUP42CrmnTQD1ZWK4vvnJdKZtci+l25PW6iUJKaY8q6Td5ksn9c7egUVYwPsLXBSTMTl2A2pqUc+5ZwK75uy5Gfc3/0rGYt9jfAd7sGMYHfeT/pVs/2kna+QHRnXUN0j0nsEfreD9O50KezH+T7nh0IeSX8t89H+VnSL/lvycQ1EteBD1LN783zDmiUZ8du+vPv/7nv/75H+/Pf9Y5DPN6qNnRXTjVeLvqVNxD0EwhuruW2VStykIovXy0J3uFFnGguoLwRQIFcPR82qVMAdD0mNm+Q+9aev9OrWnsGsnyHWc3vKmZObl9KrFQdfdbq5S90CDpnqe8XQEzGQLgqw6TwP1WzRGxOxtQYN+0PXJftXeeRqtr3SKVsNGe624PTIhu/qRzhy3efwdvRqUezverzrx5jH94LDfdqDpNeS5d4YDOMAeVa5YcRnxng14DK2++b57jGYu/0L00dxha6B+I2O5W8s3L67aHXgOvOqdZLzHdso5CGC4D0hfdoz9a83Dh7bcK7pGzgH/q6e637jU2lYUyg+kevWnJE5ftKZVItGV6BUL8+bfjPpTq7v7Xv/77n/8LdD7f8FjZz1UAAAAASUVORK5CYII="}
]}</content></body><script>
var SLIDES='<div class="slides">{0}</div>';var SLIDE_STYLE="background: {1}, {0};";var SLIDE='<div class="slide slide-{2}" style=\'{1}\'>{0}</div>';var TEXT_STYLE="color: {0}; font-family: {1}; font-size: {2}px; {3}; justify-content: {4}; text-align: {5}; font-weight: {6}";var TEXT_ITEM='<text-item class="canvas-item" style="{1}"><span>{0}</span></text-item>';var COLOR_STYLE="background: {0}; {1}";var COLOR_ITEM='<color-item class="canvas-item" style="{0}"></color-item>';var IMAGE_STYLE="background: url(data:image/{1};base64,{0}) no-repeat center; background-size: contain; {2}";var IMAGE_ITEM='<image-item class="canvas-item" style="{0}"></image-item>';var POSITION_STYLE="left: {0}px; top: {1}px; min-width: {2}px; max-width: {2}px; min-height: {3}px; max-height: {3}px;";function setAspectRatio(aspectRatio){switch(aspectRatio){case 1:SCREEN_W=1920;SCREEN_H=1440;X_OFFSET=280;Y_OFFSET=20;MAX_WIDTH=1800+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=4.8;break;case 2:SCREEN_W=1920;SCREEN_H=1080;X_OFFSET=631;Y_OFFSET=20;MAX_WIDTH=2150+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET;SLIDE_RATIO="16-9"
FONT_SCALE=3.8;break;case 3:SCREEN_W=1920;SCREEN_H=1200;X_OFFSET=540;Y_OFFSET=12;MAX_WIDTH=2065+X_OFFSET;MAX_HEIGHT=1532+Y_OFFSET
SLIDE_RATIO="16-10"
FONT_SCALE=3.9;break;case 4:SCREEN_W=1920;SCREEN_H=1280;X_OFFSET=400;Y_OFFSET=20;MAX_WIDTH=1920+X_OFFSET;MAX_HEIGHT=1350+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=4.4;break;case 5:SCREEN_W=2100;SCREEN_H=1280;X_OFFSET=210;Y_OFFSET=20;MAX_WIDTH=1920+X_OFFSET;MAX_HEIGHT=1350+Y_OFFSET;SLIDE_RATIO="4-3"
FONT_SCALE=5.2;break}}
function getPosition(item){var w_scale=SCREEN_W/MAX_WIDTH;var h_scale=SCREEN_H/MAX_HEIGHT;var x=(item.x+X_OFFSET)*w_scale;var y=(item.y+Y_OFFSET)*h_scale;var w=item.w*w_scale;var h=item.h*h_scale;return String.build(POSITION_STYLE,x,y,w,h)}
function renderSlides(file){let root_object=JSON.parse(file);let content="";for(var id in root_object.slides){setAspectRatio(root_object["aspect-ratio"]);let slide=root_object.slides[id];let slide_content="";for(var object_id in slide.items){let item=slide.items[object_id];var pos=getPosition(item);let style="";switch(item.type){case "text":let text=base64Decode(item['text-data']);let justification;let text_align="";switch(item.justification){case 0:justification="flex-start";text_align="left";break;case 1:justification="center";text_align="center";break;case 2:justification="flex-end";text_align="right";break;case 3:justification="center";text_align="justify";break}
let font_style=item["font-style"];if(font_style.indexOf("italic")!=-1){font_style=font_style.replace(" italic","")}
switch(font_style){case "black":font_style="900";break;case "extrabold":font_style="800";break;case "semibold":font_style="600";break;case "bold":font_style="700";break;case "medium":font_style="500";break;case "regular":font_style="400";break;case "extralight":font_style="300";break;case "light":font_style="200";break;case "thin":font_style="100";break}
style=String.build(TEXT_STYLE,item.color,item.font,item["font-size"]*FONT_SCALE,pos,justification,text_align,font_style);slide_content+=String.build(TEXT_ITEM,text,style);break;case "color":style=String.build(COLOR_STYLE,item.background_color,pos);slide_content+=String.build(COLOR_ITEM,style);break
case "image":style=String.build(IMAGE_STYLE,item["image-data"],item.image,pos);slide_content+=String.build(IMAGE_ITEM,style);break}}
let background_pattern=slide["background-pattern"];if(background_pattern!==""){let pattern=background_pattern.split("/");background_pattern="url(https://raw.githubusercontent.com/Philip-Scott/Spice-up/master/data/assets/patterns/"+pattern[pattern.length-1]+")"}else{background_pattern="none"}
let style=String.build(SLIDE_STYLE,slide["background-color"],background_pattern);content+=String.build(SLIDE,slide_content,style,SLIDE_RATIO);get('body').innerHTML=String.build(SLIDES,content)}}
renderSlides(get('content').innerHTML)
</script></html>
